`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
VfHl2528JlkJht2H6nrEpQiYVB2lXm2OvZhXhJZ+4wKS05RVSQ8iOxu+NJ76Mx6xIobGk72yHgC1
bHX9FwUQgg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
H9rc53tIlNFPzPpgROpzcDjCTW2aaBFPaY/llzKEwCYL4YCjHcXTG99mX3K6yIXTrAG48Eo/hCpF
bHwbjkYUOnpsidg/oQdECQBL7/IC9JnJtKwX2/MH9jEFuQzA2ZtT2uLhRCYWSEO0SdMGqBcVPyio
DpaMJ7C1zBKJhZPYVIg=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
0clNgwjN4kg9dp55JCaU5SuR52cv5l2PgSCQS5TexaPRjYgMzEwBdx6bBOtKGaNJgtu7jEEigND/
iaQ5j/bcmt16fubuZXuBu5i/pJTcNUT7H97Jg5TxmH4IxUOGBNNXClPUcpONfTGB9BCHmxHhb+cF
qDCb3hHKUCNCT6Upzfg=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
OXO3pQwTv016+zegtfnEj82Uk0jh3mAoBRcg1XOy8ri8d+x8KbP0Cx2TNtXhL8Yce6IXwd/27NET
HWTKX2D89rLRmIUWT+kFQMUe+9yxWCUvgLNyw+lNU1P4+dXORdXhaX2nb0e1G/GrIL14yLFP1pLL
h2DxRo2n/o0NW89eUJnTquyS0U/7jxUXZgVEi9ZN3lSSMrxdF0SW3r9IC86/xt6CHH6FSXwgYHFT
xG6jEdn7XNor6b0oW1ksFSA/+MxGWjBxyXzenqLqcgx2ljV6h+wzN1h/COwT4xdKo+kYbfrWhEeH
/42w6ISpNhj6OPCBwhMVT6BnU8uWr7YKowUMWw==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kur4gYBtp91j8uUNp7WNxydgn5KMJ7TrcwrpDmo2CV7ckOZiUhkAif039GukAus9f/w6mhQ5e9DU
Zo/fDeI2P8yiRg8GnM3lM9U9I1nzO85s0Hyemxu7CV17rCrEVtqhfLm7Phy171nKGj1Iiz2oWErY
2eOIJK5DZN9bni6GtZph0d6gXg+NKScOHQalaK+KxJ+m9DlowGfCXxTwVPC8NLCixFp/uYgPT/Nv
Mt/eUiEPoHrVV5eaNAohKUvD9SqCLqIAxpxT8SwMTekr4ndwFEx4eKKfNXLnDbwJpUB1U9wwKrog
LAFMiR3Pb8CsSdCBXWOkLEI1EGxfjIabX3jGZw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
jRPoPsw3+Xzml9h+N49+dhXzooTotFJae4K6gfB8drwzYONb6sN+2x+YIHO2jWrB6M9+ICj/6Fct
pyrZpFS8ViYQU5ItYwk6IQzA5HX6BKPQG2T1tlJwj16VeNGvQU1AJerulA2wp72cD6L4SIg6pIM/
Xsa8ynicAc+cxnLalQVL+Lii0PJ9Cvfk4DAngBXYpNNbQhCaU1P/tno7+DeMChrjStk1iSwvx3Yg
kJ8UBo3Dmgurg0z66qfbZsAtPZa5SLe5iBY8GlePJ/5BU3MwelNJIxEZ9RtiTVFjM8xfTx5CQ425
3yFbOmrfJhV5FBSv6pAvNnCt1fQQ7XksFK4bQQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 52672)
`protect data_block
r7/OauWfLb6Ob/S9Ldp5dtW6g9lMwI9YlUu8q1OevefxeJpucYROMkEzOI5kHLNq0rxD8EavG763
35NOLMtv4eaQjlxz7ffZrFTVqtMEmpfE5V7repbO3mGHqV2fc2+DY3rEyWC+GvHU88WXs77M7uYH
raaCly/qKsA+hWVmBeLKlQErnjtCHJ4xSPXLGdXOBF6+KbbRvl0SgQ/McsmgU1meFbOSSpuFFQnw
XnN3L5RfEo5dqBslOXYc9swkHd4Cp8Pk3epBLsO80r6YfgDYUcwLBHnOoR0yhOddcFvpzwWrBDkU
+9Iby7TU9Ba34rwU0YSz5QJsZeMNPTnUard5z3wwp/FwD7XboE55FoCZE3Cx9it+WbXMLNJrpAHy
8UDVnoGYjU2juTUhcy94f8eJ19ieNsKX2m5Lhp4kZCs48ZJk8ixHwvi6I+NKbucfSY70a5yOK1qh
Vfykwfcma52wL12YeKPt+w4RzOuf2/7Qe1v9i/ftQiHy2DPDRHtmxkHQdOqxs06zpWk4nMd3X0ff
qRA4zC+oe5REDJTlJBShtch4XdKNP7LoPyaeH3IcB4NvhvvLvnCKn6IiC6MF/jPqspvxWPxzDFQS
jTlyi5IoAotoyvlAHhKPu49NuEFYxTAK+7jfnSfqbBrcSyJLhctvPVfvAIuh8oTWLzvb8qBplav4
CFfSZ2CCEFPZk5e0ZTfrkksTm011eGHbL1nmA0RC2+zpnJqBy9O2CjZMiIWQ1FIzEUlz4eQPDG1b
VbRF+XmhCyf8GdGlOxpCTAmtQ2ohmR3/JlUvZRHtLxc3M4qGWnP8hr+9eDOvOxRobUmsJTNm1gjP
MhrbH0uoXEQVEByHPBhmZBxpoFjQU0F7zJXhNJ/53iIBU8iaClxT2sPBQoQVwXUtOl05pXjwv2ro
rFMX3/kMY7EdbcZgkqw+pOixoyHGnNhxDNBU0kSkbph0fGaV48cYTXKrCEKDz/AgJIlHsqTMx0cC
8oroIwl5ivMxEGf5wkV/JPqoMjr2p7TXIGIhsje0OPzgdFO6Q7R0Wpx1RFYcVpNw0OjKXlJXZE//
WMux+KpaMqSB3CLrPIWfI2UGZzd3ZcqYXk2FXndmMz5GJTB2XigiB2UqNUrQQTsDSQJShoNM9E/S
g0tgMM4F+Jv7kq6sfD9flcH4akeDnHAYkBVmdk9BbzOiJ3T4Z+BHvUrmRdguwFmRAg0lh9UJcAze
7ixgWo1h/cydgZ7rozJqQ17fgtXmzlmIJtEgdxvQ0Qa9/Ac0XlHKfDdWJjqHFseif2XPnCwbDQL4
OmOvuXqylobLYAt8KUyijDKWbzFm2KR6Cd0ZdYNZqPN+mVWkMEBn1lWYUCz4pkiC/smgv8EMe78M
8AxwbSVl6Ghv+GDQnalA1zNsidv/9izNno6vAhVNEfCDOeewbj1TVjzVt52aVnvB4ThJTfa40ypo
EgfdBKnaNeHsPbe7FvtNfZJ0p/kBjrMSK21UG9NDKH5uqeqwwjMNZOH4aM96+d22iscOrHRStYql
AlpuBuSz6s8T9ROijLBFexVPbrKBfwigz3xxz4IdwjQsSfymjHJKFkuGzowg/MhLIDk4NegFNEj7
+t6Zi38JihEsFbbuOAcJoSY/oEOCJov8d3zgYIxXFLBksGD2KGvLe8n0POFmMvZARCB0yYV4nPNv
BhX146riHZ+WXmdce5GVCwxmHqrVkvF6oJET6OgfzR5QoOKenPkmeacNlqJckkKGfE+D/ovPiv3B
4xIf0hqJD93DNHGMCCzG7jMazm7tzu5HYd0szN1WsHOfN+FY7Bn3sKZAz4NZq7R0KekettR1D1NO
HOLXDUSa+7KqL440SR2GHkYDePlqhQtV/679D8CttPSEhcLO2ERYN4w9lMzDmq7yobbK3+ZBqGsX
jHdKmO0o/uJ7VLiUa1y1hl+BGQ7Jadg4EghW6bxVQKRIsrWIUXkrMrvzf2r5ymc5ATRRLUps8SAJ
zywvwO453DqXmlP+/BpqueeYt+SChmxBxqGnN3fJv/MvyBi2re8D+hIAvQkgcJRGhX01qR5LL6Cg
QisZwm99O7b2IjtOph8cZrtG8u9tna2/F7GXxzmH53/QdpH/3e36UtJbHaTaJ57qSWBSFZ0r8itn
ENe+Zl8VUPJ3sqWa24tFcvro+5kaXVttjbC5I6eSNBz7SgLgzcNUE0hCMWWPtS4f/QQ3lxSZLBQV
DdT2rRj3YwbatwMZrBNhxoN3khfBID6vNnamC5NMBDztaDnYLnUxUo0+SfO6Gm5QrKWqCkvYC60u
jg2qtyR7iBxAROWg+XeJudXn3BXzpuJQgTTmTsdKJIZ0lcNNwRuSlH5Xl9njPeqrq8aTLyT1hE3l
95h6IFDi9WN7qs27QWsksB1b00OXe/0iH3Ne8UA+0We9fuJAnEqmBt5pmWT8K/SQxsM/2ZVA1LKw
Rjs0yEFWapuzgjhJ2jAPLWDrTZzZ660v8P+eDQT8uUtJMAXlzElGfHEo3cBf9iT/uGrjAaV246mC
U9N0aHTW+BcEiCP8Zy862VufHHA0gQLzKu42Yk7S90rpeGPWOpHaCPCeLbommN7Wda61iVRNKYcC
egxkfC9bZQmr1nTtk43ooyh0sH3kLtrdcTdkrA7ODGMnpiLxxWEpGsdQs88m6+OfpF1iGJOQKR6H
04zvp7qMlBpmRCk82BxcE4+pKK3AfLRE8r74Xmv/SsxM6zGqIe+M0uWGX0WMKdggiI4b58NQo0Lu
rLzLQXfK4WBKNypO0Llffw7YD3/iMQczoV0rM3DbG6HL3D4P2ciHhxudTK/THhfvSUwIKJPpKqGx
3V+k36ZuR8oxpvCjZkE8FaflZvuYj2JrY/ey7MGKWt+x06V70sXcLWD7hcXZMVAkzuLlAoztDHWx
S8ygvPXwV5KsW7sO9c3pmWFNKqt7AeqVgUl1N9Tg10gMEL2uFZywQ1FcrrjyaqCXna0d15GJojG2
gmAZC5Hjl6OdyG2jeRIPVpJ1eEv23XSnme0PQDHN9Nswt3g+7Nl1JIDmwnQTC/SNysAhClpIPAOq
Q0QYSCbqBxU3tHxHliK4CgKUaOCB6c/lraFVK3sGrjl0N1RDawheYOuGaqRcifxHVbRczHM3wgw7
1CZSZoXObL3LwutVvsw+3v1X7z60nVzwjYj0uhYq924Ln35GOELJd8xBfEY5O+gHN7MMziuQFPit
9390te9I0nVqM6oqDdlggNbhnzNmpyCtBaYj7FfzpSSmHr3A5saGxCwAU2N0j7bY1AamfjFL+NQm
a9UWGWSAM64Ljr3nn8wFa3PFBffFCVloEEwDKiW/u3y35NCQ1Up9E0Og14OgxqcuIWHVsDqTI2qE
E1iBVziNoReeed7IhQ7C6oYkmdJILLZfgnsOqqbqnT/mWVmlZP4aVsdlWV/phpg3HjewMVqBq3FO
gLdji1SnvTzOCMaYww1hydH50Igw8OHUAMpgFLMh5YSOepGqLbLLd48RgwH90JtyQmCH7B70Iz15
yGL4hsTQ8xwMr3on8ZdhQjGUkODl0vJZE74T97fawNYWiLFVA6SDG05LNSe5G318ZKKUjdpB1bH9
RIne8j9RpgcS/GKKrDaST8+8ffnXFpm/l6P/VKT/x/CC14liPEzOQo48Ld4Ii8uEqc4Mx+LO56Zk
JrnMwVqOjx8G3V/3iVcOo8tlQGu4RSW4iJKp3G04e84+sreFl3sMXM+xvaCzCox+Pnv5o9XUy9uu
lpBp/Jxi2mcHARVP8UEf6ol9ZF7hRcgYWlC54pea8gFhOcQolhzyYVja0lTSnxxdCo5bvrl49G0Y
f/hQyFrnmUgsdpfhosrlb2wVMsawvvQdXD5a7ZywnAs8r9mzucJfzBW532jN2CzfEI+Elkf2gybz
VKeT0HtEcr39CBDQj4Q0AKJ+2ZPkMW/bFltnN3bLv8Q6KkKIACJmiX3pzF6BX5AzWlvXOfzfFLRj
Rw1dW/jgl4RHPWcxFUbXrEJ0UquViMFO6q4hIlsJyIIzt9nMHa1sagjRaAlEyVFVHMTcGUrHwUUk
1bC++IAutT2aT2jXzX+IlNAOp5jRMkVSQksx6mdLSMJaM6/yUmlDF4LK8gfyrbz8T7plVbCaeY36
hmco74aFEyuDI5Czs/H6TYpI3joPh3Ppzk6N7iADveXrQL6aONFXury+EZYSUx/+AZsTqHMlOCH2
bK5Ihxq+mrwPArnsxnPnBWxWE6hnk9gZYaRAFff3fXT50QGsf9dqvbXryIzh2FwUV0ya1TBl3oQh
7fzidgqj5S2/Lk3EqYI+KQlIY3BSx1vLN/oq5ouZu2suiN381kWXME3p4fEkv7ZJKL4fs1M9NH7Z
ooEalAefMhaf8DVJEdtgl6chWGy95OUxAexPYisL8WkHTBW7YsAjPThQreWVOrAJ5AWZe9wkk3wZ
tEXJrEcZgndIvUM0la9Lloqm1rc6x3HJu3dsJqQhfcuWadh/qy1Fke3pna3pcwMbC5ylLgyPjm9A
k6UKgvlitGwGer+LV3UBbuMbuOjt6WosPJY1z6Y9J9IDye7wJe/43nr3flDHSM3hhqHhxpEF2HsV
vFmqDHa6y28byA9M9gO1hjqXVK+HLumYXupfrvXEWJH08b56HfEZAKHeq9hvdLo950R4V1u2Au4M
0ZCDJSjS+4ilKZplni3mTOMsWQ+ikxfENCFS6YGQP7p8bwdpSXCjqwAjI1RrrXFqCNmw8sq5T9uo
BXg69P2Bs6smXa0RDx0aXd01p2gDzriFpVgTSXKvJjGc+I2n6l4Vs/6fgEMG7INm+IDo9UvcOWSp
QsM3oEikKBTANEMgVvI8bTq82yo/VrdpiiuCZhCGQme08UItQ2RYCqOltpoPiVLoZhCKuMCjGlkS
jp/JxIkDdfvfuoQOCkQ6nhbRslC3htBIldghrCBxUJGtF8nZc4Gif3l4Vl4W6B0CHVxpt3qyp/HP
VKNDwg6f2FEQrFRBEuPtB2SHAqchilfLXQYRGdsFr1eeoPfC8BgRfFu9e4VUy1LZiC2Gx1ZqSrbg
/MOJ9v/qdKfUf9mONZhsKxTBpxYxe3FVnc66TviyE5HkrucDJ/8IxT2LK6LZ+qSF5y/6sSG6Yb4B
oxwQXBOYN/SeYhU6+XtXn+sOkJjWmdS4ii8JxUjp+VrQeXRowFa8pUr7rnFl0pF33xWfYBtVb0UA
sTkuDHFvwZi4xx1rsjUbHkEFA1uAahZ+lOanA3+PTwv9POIf0/Ul884Lfctbmo5uTvyRcejxVB8t
5jAR/pEcfZCsJETbCo5K7wbU9kma/qD/2nuYmqkQFZZyEMqEXs1VWhoUcXCDjKKhInPpbhRPOEYj
ALb1Jjyoi9t0munYRJNMW3Ou3hOqUPvTHBWRiFO6WG8E3me+QyIzUYmu2ZcxlCRb1StfaXlXrhKY
u78P3bZjhnOVHrvrXdGbFvaCTyxGMZxnbCattVFEgI7r+4hR+6VMg+ETxM7L+7lCOmnaPP2Gav2e
FnUkBDOgMDSbDfrhMkOY8piDsTUrm23EGCoc6MGhal8vLzG56FJdrm7J/mZBQexjFHklUqo9cPAz
/HOsG40xLHLjn45Sua7zMhS9cBfCkwWSEaxQ3+7gzXo4uRu5OUDUsynsnwKJrTF+ebqGh88mAtRd
0WJW4d+GidxKI5gZVjInzu8aGc5qY1pyD3mVASwn86PEulZYyxYB4c7Vt1tbYIerlRS324ObDdFH
/9ndTibwLsXZcPYvgOoH0loumtAHFPvxh4Tmpz73Le/ls41YAnI4l5v1/+ha8PPA80oO/8U61vxG
I3bGAowcCNpn3O1+Tu1qZSzk1aj3guTnYnRRxCXZPydijgAXsoGy2bZwKZ0u07TTp37EIkwNknVX
YYiwaUA1rHajZ/lmG6pDpKOktgo/9iKFJK2GpX+iwA75AXb9iWz+pt9IsCWQ+daGHFIWTyVUfVtr
FsZ/EI6UIk41dQmC4QCwoKgB251wyaqiEVElppLxqkfSYJ9rRj9md4cZ3OKqqLJ1zlJ6Sq+C5ger
7hP5lpsIPDECtPWAvzes9D3sKaWdLO3YsfyVDjsk3QvtW+3/m1ABU8kkLYicSOM+qm/7TWes3vxt
IZqKdjJfQg2U4csLnhNGW8PfySIjJc2MGT0Ip0GFRoTTGiyU4A4B5l3SwBiPjJ4l8hweMXYBN1y+
1QxTeYoc7qNjwUxYUWQf1hCHHupktpfFVUjkQugUYA++N/aYbiL0a5yUnhsQBoY7L2ThBJIrLRaM
jg+Zconi05h3N/Ln1FYCXCmqgqnryqjbPe6chZLd/k2OrKqKo93bv5IcoBCxHoLwjHYM222GB4nJ
Q0iuTzaYow6tvwYzwgy1p4KraQB1aZIqPVFQkXeU5jUz4WhYSS2ao+DDjWUDIpBcwStCAh0jCII7
n1wvv2Ls9uao8VxRqghQSrn8CgJAeXUIZRutg/YIdByFL9lCKFuOnCOxRMPRpCKqyjrLfkmswq49
sLwze26pkzgEDSt3WdeSNdQheRb6pGmt7BwZR8Tto/jKJKAABqEFy2VrV7YwATolViLackl34smV
T9SbEOvwDcJ3TT/yb8PQYksKmjJONhxmLRcTM0jeHcBDIs0Dzy/q4mQaZ5iWqIqMkNdPXhq7IkBK
lJJpU3tBzrt3mZz34XpDZh/78S3OjQXOlwA1ghIAxLPnJU56/pC3ENUNtJWoRpFVlW5nkaaKO13a
Ds8v1oujxpeBmzUydnR7tCyjSVJIbNRd7+RrBNIGsN6k3+mdfCIaJwBhTy/xxFWrF7StLmnhmz1d
0rWibTCxs9ViDIqTW52NBxSVqs3z+KnVUjH//b0lqUqokg9+vqehlvNCPPa42OJ7zkHdA9OI+KPO
7NgIh+C1zfJYaRiP2BC4G59rNJ/Db1KVMQAPI3W3YctbLfef/evr9T49d/w5cIuafC1TVS7w68qG
8+ZFo2oN+6VirJ/rfXvLhc7hGFRA9uxu1Z1Ql+dagOeKI07RIA5zJyuQ7xgkGgft8dJzUD/GCrC+
2CKUrpEWn4/8w4jMIXxDZEuQTWk1utC1Sg//dltgmi6QWTD/AP7CoOZVXlQGcWfb5QzfcoOpXUBL
61ahnujexG8Y92yYXPfpEK/VFKyaByj5n+nYwCHZ1SQqwd4t7sadTUr8tW1px5JSRuDJX93TOy5c
+FYDjTIKmxffH1eh1Oa7Yh0BTuDBhNkCirrB9QZr1hFCzA5frjkt5+CbI4RPkEBQ2e9Iso4aMl9h
5ddMfaJgeyT0dT2iUm5O3fCPRPQJtXKEWKq/uuldbOainYSGn5Cc4dUdi8dTubByxRxDYgbkwK9y
/RNVCFttbwak8JEBJDpxiQWOaNe7BoFuTd4mBIKsUBytJN3z2LmbpujQ0kiKwTt5bc76RXd5Ehgt
6pQYaNPJvwca6rs9MNyS8X8fQ+SESTWqbTPRyFP2qcfDlPfJSFi2Zh1JX7lcbYDsuZY7176y7Xmw
uN3us2p8sFaHPHEF+T0dQL+EkftsYNwwjx8IXc7IvoGQXL1P4ExDbkf2mj+R6gyzchfSxPwYPfZc
8ieBudyL2j21Uei5j10FF2C3bHD3fkrRWJPm6drKfc9GKCx2LoUbPOPq4KQJ3eFKLC25VG3dyuda
RuMzY/KZfDw7OvyVzABEfUJHqQ6H8/l2i/T4/XZbxW4ZUATcupJ7ClBeDM0JgQElZ/D5LARx72+M
iSU9nyIaRw1VXc91ttSJhLarF9+1bkTghqBroG0Pg101v+mbEDKdRSmGagaTuUmA/Y6UihmKJuFU
8L9iPJstNjwvYmnQhZs+JZRwynwzHXvC2rjwkXqrUifmcR/aAe+gX/yA1+hlTaBUG+WptAUYiM75
L965hApdGngPxS2CMxqMkrwXe4sr0RTLCWJaGLtmJKR0JszD+kmMPBlZkX6hHJC1H7SBEvvQ+LSa
V3H0bL/QkjkXY14w8SE60BLSYSNRutKPZ14xRTJf6axTNradry4MoyjXI///KPGVJ+ES+NgTSwNB
n4Y1E9EXjG7XRASeRN0Zyn49NA0vDXrVU4ldGUdzi5uAJWY+iwjV4yjamOdWRjHbLMMGVPdts4AX
PF/h6q/quNS2IYiYgCLt+UnjVocb0yz5EjhT7fbGFdGpVqOPVAflDkgmOKBcC4j/NhIzj8QHxJNS
R85BVkxzpLyrEiG/Gdk/0ymJigxLwgYZx/UzQWBgQRXQkprxus7Vv/++/pXHvqt+vD8OaMv++uSv
jheuPCBLsy7qumuxO2U6hPz5eUnTcywZ3EitSwXyuUM8Bc9fO4a15wYf6si2Me1AojeV4sPGRnJE
5vkKXnOJNGM/h5HN9wEOZj7V1xSWJ41X8AJ9DVEL2g+Lu3AiKqsftSdVfKSoxWwD2YuS6zGxzRu9
+1Ihm4tc8Vje4c8BcCcr4DpPjIbA1zPQomNJ7TI7ZsFyzyhRZ1C+byWTv4G6m7fBuKHSMFFIAtxI
NCENgP0s1bgqlGYRr66SvFcTL4XMSnDFIWcQTyb8COkh/MDf4oqIy+wlp6JMBniq9hJixGkrZJvK
SOb55yoLue6OdZejdoh2SfCz5+Afh3EdD+QT4S94MaC11ROCU6vok7Frck5gB2IHl3cH0vgcAu1P
vAYBzBE2vEudhdUZMO55FLDAIV9tR1/K0DDBla+w5A5MMsM2ghNGyVWqol/dxpmYVZmpIhy52ZX2
QqdCSTykW7HqKP9RNAUQXUxE8Gf0bp9w9L44R2cvq8lshJKWlvOB+0qdJ1ZJenu24KNI8gdECtIX
SRCNj+LwF19PJ7zOtMairqyIPtikPe/mg7OvU4WYjjoBG7c5Uzi9LARUJ4308kim+83636jqTfj/
/cUAlkh5pPsFwUBEBrDcvZz+YisgjHjk+VflMQ7scQkcVX/luDB7c0Zt7ZsoWYhcHMVzI+FYTRJZ
cTuelq1E0DNz1MzUfRMWqdnm5S7K5eR+3R4BDPGtB514m2d3milmRG+4L8J6pxT93c+P89fMBoCL
RFn8WxweKFO2JeVSLg4TCegQmAwvC4W4/ZgAgSKlfuawnypd0kWHmmwrAWqkKfpbTyqydKd8nsTc
dQton0yrOOAKkkE1mCUAhivLwzfLvbwVnI+0yPd/wjTlOV1jF24P3Ds6gpiSpuFp0xZhu9JPSNkW
Uvji5Oid2bkBT9xGGMPl4smDLurGfMnBhU0N05Q9gy/I8o3z7ytb/6Amf3IEOZxT2d62cQOZkx/s
8wkuVOgNMtV4sNJgTmdppiyyVoTPGGXKvWvh4x9iw1huT6tlxnO5QVETuLOk+G5lcTk5oA9sPlV3
xgbGNZtwGPSHPf9ali+YlpY3jtiuXCJjBIBHRT1gfk6Bno6We1qeJ6XYlLIU5YFfFtbaeXLdgVj1
rNfDHCvizF5onx5ewYNmIbh8jpSAggN/ArEniPOCC57m0OFzOQGBeNMwQbpdrLlVPQJqB4b6MZEc
nkOVZbGJn+L+Le5suxDH2h1WfF8vCb2YFRJqx9GE9k2dUlIpZGZtlSVFEw0hOdwzmTf5G+d/gZgO
4HAa9+me7lCNea59CyIN+L49qCeIlT9MHJk0k56w8Axhd5QxgmabaLu3kcKUAY7Wlyau+BsAjf6g
AWWEYbKwaIZmekMFPUQ9DoR4KcnjlF336IztdZcHGTax03M+VWmY4AxsWdABh6KtQMdpDch2Mxbj
8HAwxa92EA2wb2S6NxBis1SJZiJcW4r5FiBJV/puogJQlCMdESjuFC0SGpc130UlbmGtODKW914v
bbdQVMck7l6G1AZBsCfxZZkpWTMvhYQNLwunM4BqrBQwKicU9+XllYbQQsNStvcAlJGDU7yag4kB
V3ria2Yby+q2WuHIMW/ujeRdiAuVwVx8rGSXT7qJj2J+FjPqtnoAtTAKJICoPwl0pgJRdPD49MOV
PUG3wm8YwWXjnjyGAjaexYzZILCjMti5JHKqtGz0ygJUviB+R6VJu0Ifj2TIKU9CYKO8zKMxCHCx
A5To73I55Ji0nFzpfb6hm8e8+FVLWqOvuEFz7XZ4a+ZPb2MydxGmoK7zKIZKIdpLD15bTiUNUAiG
nf1mir5whSfIyjzisz+Bo21IcxoP6EfWCCAVv8DffCnidZNe6Vj7wrYbPpMfy+44/CSn/+FF6k/T
QFFsqpbkDP0eL5nQNzfnZKhMQi/aV76xzUcWpaX4Q4KQoOgZXbz6UpTQqdC2m2AXyCwkxz59EW/0
0kvCaDxKXP/J9l3eRVBqavvlTtP1dwZFjp6j3gRNZMaN9OJB0CsCYEJrN99ymG78a5GM+qazNHmC
Sjlr3ZoWl3txvlfRLOkrwygEU0B5BN1GHAR7TxVfa3seND8OtTz+GJYizF72DYlke1NdtAkr2sdo
qc6CDv66GFy1LjlqRg8e6CyKtB3If7EKdf+OE2oCy/XH9//wFTR9CwgANVdGj2ijZv2eWNvc7f34
JihzsdZoSAKzjKldLalhEUIPmYGYKpTUrjbx+iYCQJkYils46wd3zOBYK6GNK86rspuO1Gwj6mef
oWT00bPwcBypUCVzcm6MeOeH0CcrP+wHj9YmPSYuVXInx8DMtcJ1rdR86rCdwWSlguD6OQZGmM1e
y4AcpWqzXHsGYp8Ihn5XcMdoEX0G3/VFVA0u/6D2VD6X2gy0fD4p+f5HW0xJSNAbOHURgfvWRMJ8
8+9TOf/W8EsnamHE1NAiJHWpfFBdNS2/EUBJXLzeBAY62m264d/2iKNDRGiaCVUbbIj3sDBkuGWj
mLWKqGY02RYC/drt06zcXWLHXKnO+Tvag3H1IQ51NrzvusU8KtxJaGKy3a1O8v8eIEp/vCU8C0Mw
jyH2ilD7I+1IvBgSlDDdw3d93DMrS5XszFDdRDZnE77xcj3dE1wDk0gJfpKWC9lkqv0qNyxczk/F
pLJ86fJ5VjuWtyxYJBVhXm/Sfm3hqjJw1twpOE8L7U2Md2hZurG4aCo4Nan/LCJWfVCs4qIZPWkt
0KB1Xlo/2j0ESudr3nEHxAjzzMZclnvT6ue5qB90pEphkvE+h5hZ/9QGrBX7/6mECiKt8xYjxL7r
y/1VvzP0VnwHl9g6G/ARm1VmS0EFKVxtQxm0ROVZ7ZvBIHtx5/cfUrJbujthnoqB/xvYKoASclUd
pYq82tyLFDo61JmGfnHK50TUviW/kuZN7bc1WBS7YtZxJlT70+Ip1TfNvnqrdBs0bwrRg4WkwFYY
zXPjsLGinmScVtL8QXYKJ1qTxkRcCsc9oZhIW/j9NMf1088omubMWWRJ5sF/EoSAnn048mieAEUw
389NvPkLsC7Pugh29IdIyfjwRlpvv9YUAJnvSuke9N0yI8wCJ3hb2woA4snz154fY05T/XRia7KQ
LkXrKjniq2GyiEVeZ4yG1ZxJWsHFgaqlzGTknIZ2Sk9m3Kn5Gqgqt/lijX/rgGtI0CL6Tmyf7fAX
sIbnMHrhNL1Sm79RozHy+L+mgmEpfyBioJ98y4ZNmHEhnGg7TRTvtt2Dhd9QE88gU7MWrZ+ENR6V
Lw5JagguvpHR23vwi5D72QWCgXzsiTV+xpVPzRC390+Njw4Wte3MMFjNQjWm3+O8BRmBfLCGNosn
SesE5mkEqrXdURRs6hFBibWrrIY9fVVLRT4TEMzdFmQQkWxRr4vdzZubW2EAIOhrMTi0DeS4ubi7
EJBqjMVEkH+TjxdGv89aiglQWd7TCnm8040laaebBG9HTSPfLst+u5/yqvkpOCq4FujhaLlddevJ
/FVhMs7YKlZmLZFZFdW1iDzqsgcHc0yqlcLyTujWVZbnlBDNbHPq3fY+SH472HQtUXEvLdFqnI/W
TBrMTZU3oyYrMw5xS6CR+aRI2iLSBfTs7yQI/WNvn93i1C7lzIDzyOPTGCd/8dOev/0CpzFkQz2k
hF5kyjM9w6yVd/HGvVqdaT8bfRLE1uSXZXRUxyEGsuHpqVEsyPwzVgcXvTAkg8qobmxmSuVHhOJV
u+XVDZWaVN2kAugkn8KRbDu54UXYidIVnaDn/560ic02InYkqRKugJn7mCeBtnGrGnpQQsj/cdjp
hRmxTXauwt6kZxi+qtYh6rFQKd2h5Si49R22BXFTwuuPyD7Mx3QPE4PHkBWbb4d09++yXNDJaWPr
c9LTedyupknXmHE4au8Rmr9DB10+stnh47XmlIVCnkrEHlC2aJuZ5+RNC7PoI38S5265XO4g6oD9
ZZZW0Ai+KPBmROOEt/CRQ0N+Xqe0dgHiNj2FzqK94z3N+E9iTLMUggLhja4wbAy6i4JQJbpLG397
hYvibBmHnRZ+Iy/5XVaM0K29WbkKHJ5MnfkdVcMB7IlI+Fef8P8I4Ls62PPNr1X/9JqWITFhWv3N
rsr25cpS4eCsRUmixw9ZWdLDFRakhHKgHjiK2apVKpM2GcidTHGCjNYvgSZ4HLQH/f3XMq6cLyRc
qRw+Yul5aF7RiZir4RLiPAXx0BaDO8aevY68p6jukjPLsFnpVcrOaYtDj9coQ+Ak+Kb9JopSRTXq
9rjJBjd4QuV1Csqz+3TbN8YyJG1ip3v1D2zyapSX9dDmvFee1HVz+PXBMxlxVk5ieEf8LRw8KtpC
6/Mkz5zE3VKvn9FXuWTpmb7HGJXlz9ub/wo/KD/T+Y9wYupQiG/Q5Syv9gRf0KO7ApawXP9gcaEQ
xKImrpcAkOqJV8vsO7VNnSyGOpg6WntP81wV/6nzJq+mvqKybq+q4S1/U6x5/IokMdTcDfrHMiwH
/VKYCNIoEbq+dCMT+ydWisRWX1CfCNuZEC5lOQmE8gm6Bpvxe3GfZuQxm8bwR7J4DlYeNLMai3Yi
O/kzgSA9jMkHKqGasJaCJuLYeNKQg1nDna9lse1NrCFvjACWSrHGrp8yf3omTeEoun+ZngJWebpU
zXjOXNuJPs4RoeUucCgg9ciNC3gBr0icF4awbUyNRr6rxUTrE2rWhpZsBEJLW7DdrpwhbkaSwxk1
7dpuDf/dhW8yE2xRfQHf8uJArNx5nbRVYH0D8jtLdAHb/4Z0T6OIoy464OVopHiQ5AP2b8KA0pT5
kSQoU6hS6CRdEO5d8vuM4m7qArKHn8WvlUqsCb3wmtHpu5Hkg/eaXrLsbXmyoivPd8ySlzONappH
1sIwnoc+K92gFyxhtrgLN0frZfwRbAdS3AwuhJV6oA1/6iv1DsZ8ZebQH72Xzz/2u4VXtT8W39Vb
fqYazwVe2i82DCqOcVy9EKXQXPspQMdR/xXa1uEtW4oXbcMB9/ecmYPOLDa2ly1ZP2R2buFSZrdK
eccmmalHJuUfl99AQhQ7GnXnmk3qrTz+D6bY1lB1fFgCLx1OIwxx5ZHb6Ul+KoZ0TduAkxPGj8eu
9kavtnnbOSp3To6j7XGerukI4q53XfVVYBiEZnPy7tQ4uUO/ULujqF9ce8oIoFwLLcAQeY4o5ChA
x4qFtoouVt/bU+2hlhXiX99bPbEg626kaI1w9K4or16rJcwRLz24QIXchsy8qL725PGHd+KcGI/a
50xfgbkkNrLIR7stc7MVZdEm86Ktoo7mz//ydlRacabnJmFHSzoTFpCdnv+e7oUCv75ACoX0Veo9
wK1x4zRkWbljiqVtDp0uTo95MIhZgmyX2MWqQkJ0/l6HAELAO4D1g48STy6IrMe1j4BEky52utRa
5bBpFJKwKJ27lsiCNVJvCogbV1+x8PS+qM/0wGbqpr34r8Dz2crBbe1cNejjmGCSG/CN7NTLM0UW
1PefSQeBv6VxxSYqyBgfBGb05dupDSEwSM0wrYBmcwmGucgcWv6k/9kGLC6gwqFAlDMtPQZRdSGs
gcvF0hzEEN+rS/TJWHoS8g6TKsp825yO6x/KVDmi+uZ5cf/Ld3ExdpaJUNIe+TeMiV0jXh6PD5Xp
XsbzFWy2tmpGCE81zizQg/vVsUqmG9qXFDbOp3l31fdknmgA15c6lBaApLwyHVCiHR9XcNr/mscJ
G1fY0f8MRGbTq4AypYe9bYxO9+AlrTeP+2kcg4kRbOqgv9Yu32kvsgxziaa0FSVE2cwWDbfEU17Z
VnpcFIr+aXvN39Nvd/4nOQHiAnQ08HFKE0rG0kSO/m8NOk0mQkk4CpcJkfeVvIG47+YeeM6ekpmD
pnpuUUo+tl/E2p1t3U3hmifdLUVqXvEaJcC41NrsIn5OT/w2nZg122P7ALB3JGTniUqiOjB3eZ0w
uV79NchYhNxP6Fftp7eAZwC4JLgriUnRSYlNjAIMp2fRNyR+fUCUKH8RBvNRcvFCIR1XyGMPBUsU
bkXv2/sGLLROED9LNCWmJE2UiRqeH7ZlXNcU2J0zh6yPn7Lc6FecX7L27+nRTTk++1kfvLANC4V9
x7iMLqPAGUMuxlU6vEtRfR4Iq545yiSH3Jj1ucAsL5U9b8ohW1wOfFciVKvdWnf34tSmxRMkU1do
9c2Iy9NszqOjQzrzqHop8bTcjan6/KXw/qLf68vqiv2h0J/O5G1aaPphgX8QYjp+qfNqKMBhy46i
Jlbo4rLqVCAlGc3T4FNobZ5HfiQ9AVYgGljbWLjmSFa0cxr2J8/1wWlk2Re8gMpW4zhL9Od97s+n
21O2WGvwI9AvV+ODQK9PokOdUcUybAYWX/oqvR+lyzYu+pL5LBnbjtkKuMZl0VZ0Td/LuMl1jsEE
C4ItaewkDwH4GL4YfrwDjjNeugIzPDCwViCJOfeeC7P+1yoIuthPsDlID1QVR0gBsFXb1Ija/cXn
Wl8sVEs2ar8CboTtPENMTpZ5+4Pze1RTO9nClWNcKspXLTAaT8wMjtcqiu17OU7uvkWl5Kr0t1F7
s9DDT9MLTjFFyFjm8nRsC4+b5I4f2EwBvq+9wRGWN7UYjAFb1LTnkE8o+zMPB+BiYVpJtSvvRtek
i6ZuaJtiIObxr27HwcLViJo0HsJb0Hreoj+pHG1PlS4QrZYy0NPaV+rOusWMwEgYa2znwufBx4jw
EeP5F0BysDZdytD+Jof2A4dNcqfvLdYQHurFAhkwos/dYW7htidflE53OWrVw6/dEVP1Z1hlMmQD
mzyaHDvtgOil2OxJK3nwpcGv0C1WaKs50DnId2N6sEhJ84U8sVibLbvSeDCKNv15keFVKSbxxfpJ
8Rs06wxmTNA2whjdce+aHCJnaHy6mzGQt+sSGju7enFX1ZUHeLd9mWjK8TpAe1J7rrUxd2lXSp7x
QZVJylFkUBn3SjoXy3kTdT4g25O08c4YatCNXFroACyaKUhCTmVnMKCgtRhwslMpdH7GvXjB02W2
YLYjuEHaxz4vFD0JfrOsMoeLn7cVjh8dvLpYjNgt7tcDAAopi6mHUqOzcf2pVZzQ4TLW2PNNzYko
wOjcue0nePWdHVVVy4hNLQlZ1HnDzn2hp+hTHj7WT6M6pJSgRHebWrQX7LdF7efKLNmUftptvCFZ
fZYs0OR1Ywt5BugQMFpfvJ97qjOdLqeQHuSZp9FvKBl2bcHJ0eYznYHg4FZiQWGEH1L3BsTzvq1C
Fwpuvp2zpf/LWb1kf0DGRNs1NQlG76xbwdKKHu4p8oAxs06xEYzbA+O7uFkqWWOTFFsrBNAtDrWn
Bh6QBwuAUuGExINg0cM+xi6aRj0KtsRxH5QRUbodC8IMiUJk5DegwkBs+yI9yAyMTiwLUW08Dljf
jkKFaGCuUXFRBqng+pySZUlt/cX+uha8nsOE+Jv7A9B/Gv1jhmeNiz5qJ37PzS3nZqXliFIOPDO7
JudMZhkmMFFCnLPztKfr34e1VtMVi2+LpjEEmsqUBops1qtIk6r+zJafmeaWnCQaH7/1u0OCjXrT
DbJ/RDqrRb4QcPaPmuOlKGmAXZP+yHiZYM4k8nai6GL+2ZJllx88iaG5eDz6qgWXLzDeoB724h7F
XFPyfYuG1uYGd6rKdvB/3zQ3M7Pa5+Uhu/TWdPHBrrfofN5+RL6/kNVJTW1dyoAiv+I+ApJ30KmS
HTX5R7MFlBuZIzqm7Bit787oIWwv+R7Yf4udn2EU6Ey1mUADuQ+HJCz2eoDhT0UTvhFLzeh2nADZ
vx15NJa1EppVimSQ9l45bKP7OiMCRVW0xVwp5PS3ggBo63AG02BAEuxstJL8prsypmceQECk+Fks
whPyB8dlgMRtOo14TUvxBnKlcqY6HjibflPyrPc1wZJ+/1ZwELh6sEsTiq4BSyrzdiJ3O2r6S//m
XKCxAqUx3oLGaGcERu+C4qUuJ5OtnIlWPV8avb+ggODOomMJgstRnhbh5CDwOW3tbhD6/Ba/mSiy
PbZoUa70qJTOd6pXzb6sTtdHUDXjyoXry5+tgWPYiItMjYC8EM2VEQTpo1UPpgNv9mGawSQ/hosD
+66bE6YzpIi/8eUSUXefT4xjd823j2kzsp/GenrivmBm096ag3b6ivwlDMoLvyqiAsaZQJMedEfM
6nXPk2yuC6mDBVYZjXq+zrHbGbN7tfGd38ejDc4NJnn3tbCX34ecQOd3/MBi6kPrxNM6dORL91Yh
9djZYw8HAkGcghTd4xYDohH/VrxLgDbfpJyf6a1OPj++xowC1UfnJVxdTAkLRDctH5YzCFSQ5EOp
kTbqCqHh9hWAZM58EqgzpwwYcz4jBMCef7p6UcGtxzfQErLAg0RfEB07gENKTj9xIdtmlzI5G4FD
PAarCy5yNViqgVz2B2V2cLIhoMpcRmHAQy1I/Th2T4B/SeKbeW2u0+Ycmu2v41OpnzPnjSDrT1Eh
riFWd/qUjYt9m9Nt0mouyT/EofSI9+tgXki2NQV15xKxdKuhzcguBUMxpcsWCCzelpiMkRMyybzr
VL6pEOv+sb3GTD5M/piUaAuAebgIETSjo+3ycxbXM2T/aZqhG//PS25KDUlnZRRTCk940nYjjFqB
itSn6LB4P6E8hg2Mscihx0UVrHG5d+ACJah3ZrVU5xNvN5yEjxXHlrDc/jKLHAMxGYHYjQyBqkcR
e/CoNeJmzBEemgTQ2/ERs8dnqv4mVnw9fov6S3ily6s+a20ityoLRYsRxl+JULITgccelWUXzJl7
dZ/IxvywGopBsfSAGcOnqU8ibsrXKfX+X/Gd5eCK+8dU4N2Nvm2U85XDBlr3W0pSW4Eiw/JK8gqZ
ZOuP8BWaeA2nOqh7GcCCqrTHU64J2vZ/KS3t8n4QpGPmC9L7tdphdZIOeTXRas/r2s4KU+38IZ4n
TMrX8WN+89ah21TR/vTcP0OiDnRY/7+YvwbS5jYrE5aLwXxZ6ShjboJ75XSgWwiAuBISJpZjuxaT
3hUDKePwn/gehEF55Xx1NZ1eetl1CwB1J8JnOOPuONbvHlOEYlb1SXHoEHBJHzmlaHhniy4WSDPJ
WNYrPMTtXTqmed//covB1HKbp0p5i6VlaYi1iXf6KrBS9KuHTIllbRqgOSh4rZ5enoR16stzMmhV
o3U5NiL0esYkTgozc+gTgkDGGSPiRsV9xdWwOgmDqkOxGz9gNnrYaqim/FcSvusqD9jjWB330umJ
4pf3Pq2aJfXozJh96jHS5GRgD5yCWt+Li2+AC3a4xrs84byr+fn0YdURIP7qqnk9vFtLjT+lzgLd
51CLK7nFLEEZ5kzYyx4ovjIDutZnhM0tIk5wJ2TToZPiDO6cEfYgcWUKZxhhT6P6dybSV22FDexf
FtPCcY9ogh5B/zhFswZUSI7569L31RSUlotkEQIvIJE7uN24ki6gdLhTjXGJUoC4Gx/LLSPAr6PR
MWB5vswHZUTl21tsitAsIAFvAlX5ceTIMfPltenM7dBvpC3srUbqGhkq9mps8Ohx1mgWx3+d8ut7
NMYVMzETfJhJg2EYnbq1eCk0tfeUjuc7X8b5gGBMO0KjGeux31IznPttzDnxyVP/YbDYY+ZccPVu
tqQZsQVD3LGWE8R9SHXSeAiMHLviQsAkCsWixUOGcjB7zOXg7mRtE94Swqihl+Qot6D2zO10ZOZV
fycIbksYqiQktOiIGSyVlgffJ1pDNUuDiicnjEpVM22DIPSSlZ9/YQPdPIGR6gtlwtJOQDfgcG2G
V/OjTQNfMpZH1ACkQous7J1s5VFhd5uXiJbAXEetRnjvzc4v5nXBsuyQqFwahDclvWEU/eBgeXJW
H/OgUe5XDZbdqMB34+/Hv7MggTFIX7N+TeZQrvr6A4pISIuOpDNrMQYHyAK1UmtPtYl/xP7oR7zt
iGd5gNZsNg9OWVVSOTRZiZCJFDnFt7tMe2M5v/vikS10m02xJaHSTY82plikVSPhs0JcM0Q80Z/7
OInl5TE0gtt6GONLs8uH2Ws5kWcVufhvuWxn1d/TsD30PA/nBpp4rC0liLSRsAa7lxd7bICL2thn
6UfmTaG/cysQF/ZQ4n+0YFuNmiDW/8K6xpMVjZoM3mkfIrGxrIcCgn1Dx9qG1rOQeUEAQ+BgEJTf
CVsNsV3zcRpBLVNrRmyHB+htgNy4XM7yG++8aESpSjKM/nuevafsay2MH4q0AvAFKBY1PoCM3juE
c/m6M+wq08D3HCyTr0mDb3BoWrA+RnOYum7H6Deo2nVfDJmxZ4vUCDMPZSsNP4vWnoazNBK3PzU5
zRXIlxdl2Ram3Y6vSsMNBMgxkDYFw3ayIo/iYnvuYehGGKDP6LEc6hoLTxA774dfaI8eI9qjP5f6
cOozBKOTz0/qnFSkRHfMu1GTPPVtUlJ3uAOhDtkonTemgEZMBZGGHOZ9mkzL08pWJAMY7j3iHrgz
r9qVehaXjPHfpah+0BcgF9IFKGdEgdntL2fjHCj2da0n0MPUGm6clc4e8hrAnKADoqk0/zpORfw7
MCDAGxTrWr11yJHm+tCNCLLllOCNcSZAdYmachCe2GRsu3GDIg403GBMimwkx2utA+jWgjyVTmbX
pH4/xFQnayiXEkFtCuLOkDP+Ps23aKGKzV42JNIgfkSILehUVuWPYnEXNrQ0+n452Z5dp3sq84VD
WB9sMIbeoIG/SQf/aX9/SymMOsBdmzTYa3GczDBh8JFHhvmt+8i/HTVICi1lQ2wrSmvtsgWNt/Zw
VtGZXeqqLDDn/dHrZmWDCjyPvrw8UX8GwY1KNkUnWZgykrTmYQ/Zy9oBtgYJQAAHZGDB1R5O+j99
nFx9lqP+HRJhoJhjXc9pvKC8VlRzheDuvx+w/LrXam4Kl3DPUdJqlFw9bEJHUpanNDMTkvNU2qOG
qMzlLfCpV9qyQBiZdNrT8KgiBiYKdP6mz/pvNvH2k30W7YPciNabkruEVs9PUnN7XhBjSFlvRGU0
R+oPaT5I1SnOvaFCjbXtc5JrJGhL7bJhJ6/xqM/sBJNPw3NJRqFCw1W/x8aMbppBI8WNt7gHHQj1
p+i9d6/Aa1ZLkkzj7szbyRqSJRfJnJqHZQ8xh+y07CXbLcs/LaLuf/UbP+Vnt3X6jnDtf0VKgxgN
KRUaHmEZmnxEtCSTL5/XWkTP2mpVIvqkRBw3g6CRz3omTWbrhT/S/qUgSb0HPNpEMa60vXDkEwmF
T0NMAC7AKLJN3daYj8+xAivQaBsm+12mTyx+AZS/bqyHNFSjCgkQVGzQtwqMGTPknX8pTwEyeBF3
HZe55+AwACLR0nBW5CcO5bbXMxt0A/EODND8R/932Lo+G0/iltaI9Q864qUy3JGd46IFAe8+EnNa
RvyQJa2VXTXKLp7tvCyWqRsrnIIaMK9a3xtBtbTHbVFcNwIr8uOheR63Fjze4tcChPso2+D+CnS5
Vt6Nr99/pyuHkTsv5A1JRifhEQrG1BSLkxrZcx6fnVmG5WjXoMginOsip/fgqwjZpLcIbNgOUDYw
VnpHsJ+Ju5F/RPFdtwuw/epohFb6T2fXx3Hmh1aUVyzyY+3pvmkgatojTg7np/1ADRoKKxCJK2kx
atUv/dWr/E+9JqnuJI9OVkWlbeeYWlP7vUqhCOZRiPDshGCAleWVV//GlA6sMfAxKwIO2ClG4kCh
mD1ht+C53XalpRE2EPCpwxTLBQMvwiXKXRnEXiNBZ9c+AArKpR2poy0WCk2w3lPZ8V3TuTCMJP9e
Wd1uG4qVsSHOw0Hf19KIz1bGxmijKNJJOHh42l1MgnFPUm8CjZswVOTK2zearUCAbjH81b2oLUPD
dhfSB9sFtjT2hF3KMDCkU3zoJC5aFEzNfuBSb3U0BVQ3DdR3uJ3Tmtob2QpLhuqPN1veXC1RCXkI
98+eHz7+BmJcDKVOjlMlsZkUQ9LW7utl+wm8kPPDgvAc9T8FQq3251MLf0h/LPabFB0usLEH4SSL
28Hjozxlbyw5B63KOG6SnrqQcgrUSed8eRwJHB835YAasC7QMAcdhhgB/hmPaWdreKrmkFvhcLli
Qr7KXjEfnADkFqxC9zaQjoukfutQi35r/8IimeyWNEIfteQJD8rL3PR/R48OX5VfEfvO2v8C/nw/
8GPgvtX2vdzxlIpIi5+xnPOJ4GZtx1IMwvgdbWXOpjdzBxkpbkAPkir5ROzxJkQWqG4jZMBaTyfc
RXB0Kuj0MT7YKNjvsLaz6SNP5eL9UUfisJoU7OXlgH35OBN729r9lfwxnsrb6ob71PR+xQNa1xhf
jkyT3dLoxN1qo0+msej4aM+SrtOFjt+QlSr8sAnmNQ2QsWEYSQZ2qqQNYsRZasyJlaKvb/HtSc0a
rSfDDnmbzU/ILCRltQb2I3V4+4FnoHWfVDx5lZegsBfzjRmPol6T9QjMC7SiYNK6UT0AYmEkNEN/
P/8PIGjCsL2yo84LEaazD3n2wcQrtuh1qFMbUXmn+M/UDOosSqx0tA60Itwk0E0Le/JUS7ZKBK7D
MJHyGnuuKgUFx7HerL3pc5q4Is8Fxx+kOmjXkAD1mj+r3/CNUEUALkPStkHpIcsx1jsfs9rdJUi6
TsQcQ8cnopO2LJSnHlklbnfc9r1jjaARS2xGP3bqwK2veHh7lhxKihg4yTM+TAJFU68UJSIYhVEW
BSldO5dVvUDFMLgfLthPeK5K5GCFAIaSVADz5jIVxbVk5l0Hl9s/JKNkJW5j3fjZ/LIqfKnhNHSH
NqOazCTe1M789ldq9jiI2WFOncSTXsFQ17NIG6RC4I75xHwLCGQawCAx0x617RiKzyydfQKwg9ZT
fpX7kepcuUk7X7GjBFFY5tIdBl1wd4mFA08zh5t7ywdIfxT+/SHh0gQInZSVder3203honzWeiT4
SyknH7n1JwNKMCmSNWcmB21sTP0JyieROJsOdNHT62PSirBOKI0GtohOlnCIw01Os8bUFPohyhA5
mrd2V1GZO5OH6xvbhj6OgnavepgC8aUrmxVcDISU+4Va/lTkkF8svmoQFdbhtfz9c59fy1vxd1PW
po9EaTHjnec+WA/wCLqv7y1GtYRW+EEQi3sPorRMa0JvC1bx3gseeYPtlrlDl7GVouIL3xDepZdA
8/39prUGhiSfY8dnLWpGvjumMlpExchkATXmLoqyZQ4s9Qa+GLUPCql9ksigI2bZ3+GhUUv38OF9
wIdFTezN3v/lzu1klP6CAUIRZBI9QjMoZ6ich4FrXZ2JJyy/2Lhy7NXDvmACC813VQ5mP4YUJVPh
3nFCHOG1FYZAzisiV1J2XfiPOyRDBvwjyJ8cjf9ECH5HpX+oyA7B1hN+426FfL0/NHiI7+3JVCRm
enAUDcqUi/G4wxUY5jXi25fh/RScrgkvuZRNtM76oAo3d13ocD1o5K5bo6gbLg03cpZAkGJ5Psgn
gUrM6LjPM9HwXE5lX1y9XrdeotkBLLltjBF8R3JrbDRyPQZX8wtHjjS7DuRQpEFPl8Q/Zc6j4gLN
ROxOTWGgkUmrYAXGwg7mYYdYD7B8TfxZh141wjjFssjgqYxF6EYIof+1lEqdJz+Pr2kBA3U53zj6
UQdBS+S49x0PasX1SY3DK+4GksUrE7CjPYGv0ad5PSJXFfgEKe8vWsUaDQh0AotOSK/9dizqgstr
VTzGEyHXEx1O867oJGwmAFe2fa5VjBcZI8LKBCGjajAwNwFPxAaEE9O5W5tyOpbnVS30OkMPi6mp
qtCQXzO+nhIgB91zkD5n0vog7HQAA+lRGRkhea/MzxdauXJdKVacOJtMXNRIyeK5jsRtKFs012Kn
H0DvGfBvRStc9yghVvtvRFODoqwb24nLc0aX3wzC8pkuSgSdJjnUUQeJV26EM6aQlpg61MoZr3Id
5vWXBuoy3AM5va5pMDNJx9WUyyjyNzggbn0/xc96vPDblDFKcn5Gysj5niU0u3jV3AC7jRxOo2pU
2iNmJBocXcwTbCOtZ7FiF8jgd8KhSj921T7dtuRyq73/MTLRhez7ijZcEZ9JJTKzi6gD7MITgIRm
eUQmNmJGMIa2VUALuFuHd4dlk1ZU/vixK629HSXcyd4SDxR98fIEwmDKdSs1H0BJG9ZIaCedP3LS
VLKPWgcwvBxp7jt96FUBPPk+4nxF5r+fOPfX+1ITAkrochuW18Zm6oW0svwnoa4192SiY+WIq8KS
tRqXEDzENNOOTfZ/D3wKB+JCHtmyEjYQ0y9VBNd6xWXzZdZ9jG5HUoBVdvWF+vi7aU1uJqO9RyP6
qHP7EZQLPZU2Vfp9fDlYofVmxWVxmUMb+yZnFVjZy+gB6NLHdoLl2By5QzU03UjpZpzYmFVh8Ca0
dRsnGTjRicbz5+q5Y+RtH2IwMZwj9Qq5b993H41oE5LMiTFt/fhaHRUnOkzHcPH2SifFNYKS/h77
Rul41TVmY6Szkt5huSULKBDrrx6nwGA1l6LswbdGXMvoWR9R0UpePlxxvhPekDaPn0XSYGrh3FDN
RrUAZi57/qKKu6H1HeNnCcik/8CphFgSFSz8hNcWljUWBfPIBUCZmQF10gv43hXQBWB+pp/87MSG
No4MvPgQtyZUnu2GbCbvorpjEz+fNdbaEhY3sWY9Y2uBZN/T0zC2RHDjS/B9LbDitnq4rwl+E3qj
ulaV4GOcp7zL2WSNa6EyffnYjFl+GvG5jrRji/i7fyI2uA1KS0n9uo1fkMW4QuEMF6Us/CQQCak3
SSNINm/urZP+bKffGKUrKokc/ZQkVguOjWxPcScCbdaOux6wuTj2Sl7TplFMBEfuqr8ugLAs7dd8
b2oK+C26B+pL0sAjPY9zv2XVnv90/x1rzrYZ8c1RJsJt7bl3s7ZEFEf3fBSUQI2UdkjRabIZNvaC
Xad4OUVrUXwPvFxsPFZTFg4347e5hy0ltIaDBnKkScIeLJ/vkZAxL4S1ZB1Dv4crhtrMQaJb45tI
JAmfsQpuvOfonSnIDQjCtsFnF/1WthMJa8pD3bAcR61UIsjqyLAmtT5kdq0ebMG3s6KuuIV0B+OY
KIF/FtPUR+jk00nELU0TqASVzn0iibZa6pX3tjnRvqozNBAwHHZ+0TIGdZZKb+RRx73RENyQNdza
hyJUnpPnIyLMhKKoQH8CtT6gUdhM2gk+L7mP9u7MPRzepjb8z8oqA0s0RSdX7eGBCSNsQ1rWGSYq
6kJ10LhpoG2iVuygeKQjZX2nQJeK2pyruPozrMj7ooa+Lp6+uEcb4/RbblJitYbT26xK4lIXQzHm
j/jS6Q+kKS2LYJk7ymnhg1jXY0mxbDjK57L14fE0pMTCS6e1L4vmrB5+MJPTaedpyQBAV4RmChxi
/0OAwO8ekbaN68bQb8dOVHGmwR1ZJ4uAVImfcgb7mBn7vvTWiVIE68LhxhIlw1vcUOr1hq9Z2eRk
nPtBLzkyrp7NojAJw+rGhfRzY6VcKAm6uHMwvIFCRzsS2BaA7pGmGwvWweS/XE+siazzgm3Zt5+W
xZvNd2WvKuTLrGan5YkItoRwbyT0/47WLCpAEAfOHTQV8Z+h+Y9XfWz0NGfkJC/0oA8I3Yby1LWG
WzkKMdmzGK4CZt3hwWXeBYh6n5UE8jhGVpYqc2kExEU80CjmIQoqN2WYT+S9o8D7FJR4TastleXQ
7js6gcvS6VKSFxqy7ocD+l79jPQyFjxS7W2zgwv94djsopMe1zMofKWH7t0V9ny8AIZy4+p4rO3L
sWyHYKmhzXrYvlw2IzApZvlsetqlANlGQn2H1y8FSwseLZHDox6kmZQKepjfgy92Mo5YKBipAaDc
z4n3IQFpGY1A2iD5ULubLjHoiZlMHL4EAhfHdX1BmxO+hO4fxPYm7LBjxJ6B3ZS1VQEMkKp3SHDb
nxgJFci6ECavSNcX63LJGnLFY0WmmORwqa8tyy6FuFRUuUeY2stXe/0WvExucOi3z+TOtffKGSke
yCOs1SL6kHjM93gc2r+zg5ZV3a7E6LgxLdihmpfNjZpPRo9yqto3R6+RMgn1xG5m1xvs1og2U3wM
hdFX+D23BEyljeZD3Mv0WHEzxLW5JHgP3LPOiV7dpjBwDxtD3yuN5z6KkEhL5uhdLHQNcVcFn7yA
rERS1lrmONplVOVnVSuQr4jEL59VZHf7Am/odQtZKJbSl/z4IO3jvPKGwFdhAMsOON6LbUgVAxxd
VGFHnxsCQPaVbvt3Wva3o24VZIBJ5SY7RAYlTVC0x77lrl+d+5JkfbuO3wJvbGa2OmMW7And9M3n
7jN+O9wzvMtD9TNCxf5OGQh5HI3aj+6Xb0M2CiPpkwwd27j6ycqpu/ZJOhxElKHiSIlGskIAWoqW
BSrBYBDrPwgWSG7vr8lrSO81/eMXKyPg7piL0+QewgQVz+SYcV9le+sgU/e8w8X9xz/6udir52NF
534EAsew7ui7mLrE/nBaJcaMtG1K7UBm23k87Ex8y81GxBWo2OpOX/Si+S+Gg9Me0Xvf87IXQb0U
wG+l4tJ3acpsuojBUJ99KLdkbJpP00HGzu3gExMi94wU1hlwwBFz4pzDJ9u73iUy3iVfjn9d2fZw
6mYIwqHUk73qfYOCoOYwmhQql9l7ii4FGjYHHXh4arEMvkr87xoRbx80jIApieosEm/gdB7S+OQZ
LPUjmu8aXI+UfZWi3EV0Ev1eI8biJ+DnMMOYIZqjNO+DOtHUdQqktiw2PkNPwdGmfUey+v09uQPF
mhNjkRR8Upy3dErPEsNrvGc1rUSmJZpeJcrAf5i9k6baTPtoEvgzWnBsAjI1LDut2XwuDxvbiy4A
aq6a9DtCxIYh+TFdz9ytVG4lvIJUtvI79gooqxgA3GPNQ59b1zYXlMbw5WQv6BtQd1gkfpKO5qbk
9mqdj+qAddYuLLBeJ84yZ5CuNDcrtdH1ZwvfOQTNgpdUAmfoyoDvrcZUzjk1H0svhsKWzhKPxCaZ
IYmG37GcThk15rxawUrP/Ps1289haWEwnFL0C0TEx+KcPMVtDIDi/dEP06wOO7RXbJ2J/0egnxKJ
w9jm/UYQGnayOkqFbt0yFQZgopD4Q0wlMRtt9zL7YcW1B2qzpAkh2rMgUYUzmR4XOmOFGnsPa8UP
i1nTh1bI5R5wh+y5UHG/fuAW1RdVKu1Gy0JtKxpNfxwiubaOfQoheNG71xiE+XFWhqpSImcvkPB1
15voK0tTzRqCrutfKcd2Vy5KMkNDmKBLKay0Z2TiT1GkpUHSc66dXC40SKHMiNoNjqplDabx7tEz
UAKdAT3OF2E0cF3G8VEW+FogeUhvvZoDaYtWRrzjyX8fFnz3Jz8aKdLXzSsxPR5mGLtk6uV54sq4
UUQExuTKKMI/VMBWRD5eJ5qxpSJ6Y5LSSEWpLUFU/37vNZH1mtVVTsZDNsO/QTZM9luGwZtEGDH1
+8I+F1BSSwO1L2ZngSUpffI7KmKuXv6kwbe9Tku0pAT3lChab9lBFMC67kqJUuAb1m5RLTctGAij
Km5Wr2xDlH+zgyF2DThuThJUzqABO9mx++XKoPF2Mfyt0D88/h6G+qyLs0NKFLJzd13WTZrH/8bm
yWas+Mm7EJ+kGxK5pNNeUUfYJuvih898+NQ9gB2eTJiBGGT4TWWWy+OK16ywf8NiszoWOZDZABox
o+wPY1F4+BxFOFRcRJjumErJgMNKY2YfnW3yeok/ZbfyDE+SU8BbqM9WdCsiwgpoU5E43JlwSeJv
K7rOTPs17ts/d7qZB5XcbYZVYPWGuFzr/0es8nq2OmCjkxv7n7eIiGVq/vyPfiKSamZ+g4P8d3et
n1gWr1KoEZm/ZMZMwLYFx/Fr//SdSjolRjhcqSBtnwQC8lBaQE1FcwiRfE2pdvnHN3o3o/aKi4uY
PUHDhU9EDOvnWzHOyLtmV3aR8qeXhru0gzbjT51IpfnT9OYXzLdq4piC0hHw+LdfYmooU1SAWOz8
ToauvoXJ8Aut9WL808DwbEPcFzklV9T8SRGibBvLgGhVq9OwLT708vjoGZxzKwXMme3DjWM+csAG
1XPiDrxH/7ws5+uWAF2d5/wi1plzctUu2MjFQduoj5TzgnfU1I7KabKUVWVZ0M6WIA1M0j+QTO7u
lkbnJUn12yaVpScLDZyHecmVoJavlv8Ahvaf34KnCat9+T24RMaqtr7GfZCKkNRUa5LMBnTaRwtM
rYxUHq4lBCcJoTnk8sMi0IUZBTD0vBNsyLxeQHxC3Utvcvp0Ko8kLhgIOkYMXM/QNJr/0zpR2X2s
KiKBFFu6/2bndTm+J98zlKWQCm53hxlbnqOGQ0Zlwt33UDdJdren27JaAy67VfJlNBCi6c9LQIZZ
EHe22+SL3dTxbuuLXkt7QNi/4VYRCivWaQkb25QjXcpt21JcT8LCWhnWEQ9DoZh/fOFQbgMA18xJ
WQknXqiOZymP6NXoH+zq52rm4G6pN691bIK1xhxJm6eakR5tMETr/RaKJkklzzyvT4uCHtWipaBW
//4RjGdW1tu4G6irw7YiO+B1jkmmF938G3U01uflVf6KSxPjS5LWAPbcknANjuuA4dO3QBrgzOeg
rxcslzL5TwWgRTdVMbnhaIxL2eV4wIm/Es41Woo47nvL/s6cpDYCC1DA+DD3ZUfRsXKhZPxQE/o+
IULjxmlHaJjFm8wmo8eIp5z0TvsyJ+7mzc6VhXVtmnyHVaGsjQEd3LgB92erfLpgV21TKhqBdZNn
BrQgvR9KWCEGEgwCoYEBhx8gCtbM+ASkYpFiqvalBRSCpGogJEknoy1I8/wjjPIj41YWyStwXX+v
FASM7aMdASsk2+6xrxhsZita5rN05Xv7Q7BFfewfdhIld3K1e578xn8qoXJpoecgB4GDzlqgbQ2P
/We0VeAFUFC2lBJ+/nDQCfiwkdiA1TPH4wX8XkZuao8hTUPNItS9o2oZTg+H/WSRZ3xeK661iWJB
4SMZ0P7ZNjGSegLABMXLYNZajPh1Yi1ON7YTFdCI8d3NImZ1VuLVGLuNEQIOIBrL8XJyyjdHoOKN
BEttfmTYHX3Vd+XQuMZaM4iekR+8eut4L9QQYcNJBJx7ri6W4iU3kUsFXrouJPdFgYPX4bRgeA29
C5iTTNX385iiBis8TFjpcBfJ7CEyaqVrMutg4MVLTBaNrUV9HVpH9MOu7vww+rCsZGleNUz2UjqH
DKZLsQhVjT4OvRFM6LXzqsNNQLdIgYTvelnySLeVnrXL+UPgXwihxhBUxOlYh6SsjxtbadQ8EAch
lwl9YvSmp3s3s/EshNbUdGJsnQcTCzqhr9F6ZinUFr9CGNUxeV4MkvbT6LaHEv6AQRAbHUDRFL+c
d54xjmgQz89PxnziMYLY/dTk6yoagU+w5/fs81Z5pdp7JJKTUvp3+Rwl4YHcteIzp+k3TZDXNX2X
aTMmSbuz3iW9rblKNntv7WY/PCNpD88RlMzxirbUUV29c67rnHAooTG0Oim+S8kg7mbn9I102Snz
7XpBAYcDd6P5dnFcxPPAoS8XVFVgHsnwQd0yFfhCXQYRtUwIC9mz3RaWuLS9FIfnbMsCrD39mEMH
+GnvHTs+KjMFvqt0SK3uYfmrDkZOJe8HfuKMXle9wPdYyRJM8hjF6lmFiBo6w6EeHw2mp3Vxjkt3
y2VvKI9B80l6ZsKObEln0uwEtCfkXjKKg16g6wgaPdEHtS2WOgJEt0gGS0RyIh53GMLvFzDrarZ6
Z24y5iDc2OMhCxFnZEab0qA1hQlW3/oiAMBZHGrDja3Ps+/8x0+8PXyEe9krnOGGar5L4HUedTrg
aW8qL5yCCN+4ATY6p4dW91SF6OicJvVvVslUJShka/ORBzxoHECcRJfj3kgmTuh+lU94Z4vqKDNQ
YlzZJWYskTHITKE05QzG93+2MyiAVXYAQeeKt5g/v2RSX+zVdVv+8reV3aa7JHVG02YMpKXpf1h9
qC2L11tFNmcwVqtl0TK3fEWiLP2tq5ijI4T7z1Es9R78xBBQbEDJsvhI6MonnZq/TNOjH01Iq4wR
R2rWVBCkEYdzEDzyzFFMI7jYpdYChse83D5spWst0fzuua9y43JHoG+LYbXGaGiwSwlBP1BTDR/5
0VVs/tEOi+yZlcCHDcxLYdwpDHPf5zONIRvNNNWDwfk78Zi8ixm1oRACgi4McG0pIf0orkRPEFHE
YWE7bbsGIbIWI5Tp8nc4Q4707o7ImVgixgYXdIxCm/HUJAs5oyVgkmohn6PP+pl+40ApvpGzCBVh
tuPr6GQfxx9gKppTiogDlboeUs3x5oSRQnqKxaueeHueoajw6xMHqHWxBS1fnOpyMAjAu4Phi8Yf
y+snk6IotNP5zbDX7MQ9C1FY4INygM526Mlz60kEaUWUIgOcuSiHmmdLYKwpKW5sMCC1juUC3IIw
SXjKc6lq3Ncjx1GuYlQcHu7iId9+D85ZRC3abosHmtYWZf15k+TxR5AOjiSEZrJdDgB5FtLFraan
x1v9+MfmaxDSrA8amvvd21HhPdeXUjPuWwoYYk2ibMALHRpoZWovDz7Z713wn+995ZOK2yjwlTRX
ut51vVA/MYie6jsu+BTOUWrrf0SIublCYHIMSrdOcuaZaqhV8keohzGiOF5DfctLA0nEZkYgHR3J
Z0IIwfshusyMB/kjlz14ZsQ7o3ctjqv1GLpX4hvO2kmz0N3hkqReR8jBNoXl/tfiMRQN9C160u7z
QfFzaS/BsBqeq0TCKf11CXS833CR+y0rYIA34lQV/JlqJfhphsLFMy3CUoAIPAs71OLkYHJQpv0/
yD45Y31cbHVa1nVec257Zwpw/w3JeYwlKv7Uy4kMMy6rZjaG2TowINhsoJ4tMAU9mog3dvwP6xWY
Xmo5MdUQBF9TpYM6m4GT8GIM4VEo7v1VrCeEmsa1Q/wZeed5GHkoCZR3zFq6XicqJK+KX7ZAQeWm
QGIbWAAYaSQZhvv8+pVHmJNRGseFY7Yk+2qJiBXbHEAnYFdRd3jiQEtBcRksiUPNP94Hi/PUpjil
kC/6EDOFsAdwyzQUOoJ7A5yoUMHsTCA7oxYJTo+qBgGCaSTupArv1yqKxfHX8I4EZyU6Eg445daI
sKTOdfiJoRhg2ZsYhN2eOSozGBBj1M3OYMXCyuXjCVrpYwjtvyO/y4rA0WgGZEaQ4bVNdNFeBL2U
dkvbHtg4aUGVdt5mmKckCgFkEimPREDj73G4KAwSZUHpQUR5QZCQXm4JrAs7GsslliIwAPptzlnX
zu42FPVlLrcYROLPKIRPYXzMDPjyC7quN0LBjbJnEUIaDFKTNJGYPWP8ud+jsPxI7wvrroUBM+oo
v8LIn1bTTC1xcVqcsDlSWaoWsTFWzv4RDZ3BgCLkIuyd4o+jHBe06nEj2Hq73xNVRuMtG4aA5sBx
IidhwjGyA5DCZ+tpDnQ/6neUqJGSbVxUczMyuwg+w0PQSI/hBur9qwsb8pfQhstrsNusLDMZqrT5
yPkTQaAf0i66QfHI/TG4lxuJB3BuKTSU95+LaYjtbAmFyxZbziazFe5qYL9lAS3h4go9zjw/z6ZJ
UuGxzGl4pyw0Ey+uxPwXTwBuzBbVGM83sclRX2KByAd1BLpl9TFQn5qqSXttkxGn58mo6r42Fthh
df6NBiPsByvQOV+TBVnvImEpV/hq643cQfGWyQsa14W5Et3NMqnV37PI25WtkZWbZQKxrOgOUl8k
90iJKp5L5aF1b54Q7SCMJUyDychv8NOLB8BgIBQjFNLfpnbvAu8ddo8g5e76HyHU6Gag3UH76nUy
NY9qdjcEVCm6lCe+YRGNzDWTNSOAfcT9PdFxiqoqr2JUaPm5Y9HFEkEa5xznhTLoge54fbCbwrD8
eqj7t+08ZF3UY8UD2k3BTZ6pfTmZ+iLTqYIV2seCQTeFqF9R+Zf/swefrSHqQRafZGRkAH5gehED
ZT0SWYIPEmGoy8g211Df/JiyjEEfhMm/DlrtVEkGkotrV5eO/HMHUTQHtIy5ai5Wxl8fc5f7DK/9
S6Ga89NZa38Ky+E3i9v/E2DSIHpQ/cNhULzHjH++VQeJLuPx5Hy3aya8WPCrrP0Qiy5uMStVxxQO
w9FiFq+QTH3PrxNlnwmSu85+OeqkE28kxaq/bA4yoAxw3jdCWZBRlFe+XBnB/2VbPsjkzj4HcdZa
lmu30j2OMmU26zet0yaGhU9z0zIC02CEAPUDlsoyt+HxMW+cTGpaG3kNx6vNz+s9vKq0ApFWnwK3
W3rfD7LKCEoLL6VICppKMz8E7vtpAFBxkWOSSIY5zrt3T0X0E5vtMSjkJRRi8bTinGuoysku30Hj
edeANbsJ/sh53wxCn3b5jngkqd9JkkrczOMSAf1j7cSNb/vfuwpM4njgjWMS/pKuWcpnBkibwxpC
Q2c8LuyUHiVhv98+TlJ1pSLskrk870hsvSjL0EPmWYUkvsg18Rk/NmGtkAQnxRYD8Hi3I3ckDoeB
kaVv67ZAH0ROT/UDHC65t74+9SYt/+DE3iNcagfJhRnyW/2k8uHr6IAxZ+U6P683xOxeepeF5ted
mqAG3Hs2UcOyyNX+47reOqzgknzaGOxLQ58HeJu2OegBTDuNK0YhorNVNTNQmLZOvYPD9xBc7vBx
SVf8xPDX0gMOjYzD6KQog4g/WJYpJUavk3MKguepK4ngBgZFM9OAFBFxvqQym3NFe+kyTFTD9HZ8
cKS+ZTPpwVwHU/am+oc5hjFQLTp5NPaO4MwqSqa02ztsnOxBa1It1xAE5jkKRVbyRihzRWVlxbDJ
EpMSCwYKjD9a1bltDk06HsYHOwEa+OEkCiwbLtXxkibf5va1agEuMHbgjxo3A63ZOBd7bp5QtVg5
UxJ4Qm8aexGYUVHdudbGpBmkSPUqdkW0HqMcNPB2nPkUZ9KpJZMrnd9/I6Jf97JH0PHhcH0wc/hQ
cb3WUg/VoEsj7l1PDJgI7ox21GSvKGjO41Oza3rRzybmXjGwosI2nk39aYSi5JhtcQ/XGDeouaVY
ZHeb7e8IsfdBk/z9g0OeZammBVHqL9haDVIaf2eeO3zRXVoafKUcCPq2mMRB8eajhSbmlvx29Pfo
+JuQnxUGfbP76dLaU9EZUm6Eyu9hNeCNzPXiJNu9BlgpXvVgFwIvd9v67WkiGz34BfpAtZL4NySe
mdO5BBVFypIss1d+ByOlerM339nSlrrznDNZH9578kDPwO+IsUp0cRH9VTznMAcnrsa3UjGwy2t0
JZ6qgr3IEgkmyBgaYHIdnUxooi5G8XUQW51b8O4WOP9H+iCPigJJx8WrAn4ua42x1iH2j2VVimGC
A6ZgmgIZ3/2B7NwjoZOlAEQRESYavcrGchyfSTUNl5JtYRBqpKRYMHvVL3v7GVwGY2gn1Szn37kV
lK7FlQuJWlKSiQpf4zhbfYqaX/T4qbXxOfmmGgfLCfNQoUNNWhdWcHchivjuXih0WLI2WjYp8ghR
vGsPzdDjKqcPbv2llKUqQp8yjX/Z0HYdGC/HS4Il9Z+nvy/JbMPv7HwDXYQobVNl7VEsXOfScmlF
9ZMqVvJctkJSmzbc4E4/o/4mylKqpFNqnBHVAYqOUwBZvIy13PO6gJyuCkPhwiBCrEM5EyL9TEM6
eUEjtmeXYYFh8ZKW2bY/mY2Q9e27ReJdMPquecaOCW7GvcFmtXxjbKiuwWhkJUuaxg4GHrut9WWr
MyWkNw7+2iKJtsOaVLQkcJQowXlvMchCTR898i7O5fLV77ToSTvU2R/kiw1HK1FqmqDjExJ9B8eN
rMFabpoaeGb1m4TqTrFdTvBhJ2ETUwDD+BwSJTC7gxjlvTD+0c0Lzd3F6OVibMXtcIynyTapYT83
43uKfwEEjCUTydH3vi4oVYLd6ISpgj9AUL7xOjdQReT9/LFTBdVtju7WfWq0jNHkROgs7i5jrYRt
pCP/LubKTmRMYorpqC1rUhj8GkA9BB2oCc02ZcQYB+2BIIY4renFD6cDYe50vQ8vtETVc+cafls6
WzalC8pB46l6iYBubnsfwwXTwDAfVc+wkwAPiFYW+818VvcyHr4aWJzgQ9+W5IrLTos4vQsKyzR0
Oq7n6mW5C4f+Fta9YQk0Tii6bPi3aasvUYn8Mv6IGJnw9bgfvz7jo4T82rmsJU94GQHe6U3EyhfZ
Qid6NpuZHFcJuXDyhC6ScP7RQqm3vbU4Xo/V81k1KlUxc0zwk6ELYuRLaodP2bccDZ9OdXGCgwZC
9LR3VweuhoxruPKakFx/g1RGD4tZ1uiCM07mDjgPCuoeTTRjmyzY/QbaLXtlaXrV7yabDNQ1VF92
/vd3AKW0g1YQyvFUmsx7zhH2muJrW3l93oQk+VrPJmma433g4YdgzBLbLFRVDDRssTVqJDhlJmV5
1BK7+Z8s7b4NEZj1Bd/aYGSKw3UQtbAoXJzPG2paIfe9rPy5p7OW2oy16jZn9XZ76GDYUY8lLbTf
g11dYDvxcYQY4r+vyI8tsJ7h5rnj3FYUgqH+F6UL48FalagxuXEFUmfqp/QCqcaU688Fvus9bdUj
c/Jvlh8n1PfDuODLhmgwIYDZinHxRrq35skX0NOJRsipizHyCuLRYL9dolltmMmTVMVho+px1I0Q
WcDGV7NXusoUtEn5aTfgE4ZbbkfA3IUIY/JP/4cauw7so4gBqIgTNYu0omXV95gaEmrlM/ZwpUlQ
Zy8sUpzX8iIbfncyXmoOLatv8afWdQU1Vxfk8l/LW1ZATYzTEpVeyWYrwZ6m3NV+dtqDnIKHCC5G
MSh63d1KbXgl/9ul7JWVpfwJwVPnqbaVuL+GQP/fm3s8QKdf+wjPj5jWzmRe4hXDL+8BNpcHs6tO
DxSMgQ6PHCRmgzdOMmDhF4TzjcVtPX7F8ePyQbgm5cTL4jHtrVc2mvEnWwwenN4Uhq9NvIlbwyrH
HUrXRwuXcv59TUoaDvH7podQywyMeD8DPXC3Xqr6F3gXFyHaxWgak2mMLSHtqXjvdPP4KTOfRMXd
HCGdvTryd1qbe2jpRIU9bQWioLuCAhZAcIWragzPub5Y1YMqLXSAP9164ujTcn2IMjE5z7/1CW9M
6REjC/tZyav+XDITJBxOVXvnwwXG59X6Al5qaunagmY8opo37cT5FoOzPmBRssVXwr8+frn5Mu2K
Nv6vE57gvH2CX/ZD1plZdGBx0VNqZb9WrPlBlDM39++VkQzJFDp4YxbCeUAr6PhABd8Or91L2r10
zTa+BB/lFD7tthXTgqhZEgjxO5WP4oXURiQN+5DGJI/FRNTyr8tgC7brNXWiAuzgr0u7SNvukkHn
KyIZRwc2hpWafJM0CZJsJMyJ1JwM7shdf+ZP9U/7p/GfRH4+Tv6xjGJDsFCxCaQ8eEvx/jrKf5Nx
4L5uKzm08HB9IlI+dHe1F+tw73TKf5s705/DGDJ0QHje+noXGqwUbid6kGQYBBbXaRrPx2pFuH/6
5r5qvrUwcq2gBKFPiOykzzxfWDLt0y33TrrEM2pyCvO9QGqTo4t7A2wRQeRbKUNcGH/8u6ErMlng
M9xjIQ5FmH1gV6F8+OkevbcHRfl7Fm1oqWnKiqZZd5q9LnJhHpuKT6lFh/0yOG57OyhLMgDgUPfw
w2XLGKLl06IPtqGqbBpXPC4df3duuudE2ccT2l+EPjG5mh4Z8KEJ3Kh3RUPvn75g8KGjEykcwGvB
pARXoy+9OSSBF5XL5rIy0enykU6g7k45Q47bsxYUNBzZfXsYKKylsFUkiMDnnd+7CMg2CQRMHL2/
POoDBAtgZtGkSEIfPnaHlve6fxTkH8yFj2mkz3wVAjqcZHZXL9XJDrBSfoLibq6kC19a6XAl/7Cs
G8Hoxmep1znKChzRk1fP3OKpgfXqUz5JLRgOXEFlme6s0Vg8RD8Il0l7fzp1AYIQEGl+3MiJDBho
XCaoR9ufURpdd8C9t/KK5BnCS46rXN/TUYaZgHEX7B4V+TWHIIy5sGSryhqPNktsuoOta3wpUaIf
3nz0Oty+2jmnENmRR3lLhyfLLB22vPBFfdoefrn4U5uNlLtNA0M76IS5+PFw+gHhdXXbkJ1J1BA1
lx8aEbPqMgHoF0WYiRreb6i9Fu7tRaHyx1zJrvA/vxHGP9k2nWpO+f6Hd3z/ImXx8Uh/2uaBirih
S7vXdhlkHtRatKA0fjoaM9IKW60F9tupLBEPwbIS8nFPycYouI1hXGdtW1GiMr/TeXeLaVujQbts
apW6m5wWVaDlzHqESURMKP6hdVE82nxCJ1DvJrtWraJpfFoCiN0sA+cKt6Gt7V4+V/UPb8aTt3AA
9OrZnFWHcdSXGC0LkLL1KmVXxRLZJ/b/lomUmrktDx2Dt+fFa3bT8o8uKIIuFKRffFJb0B0ZNMOf
gNhzgAZft6gzQNHp8To/S3BUfK+DU4B4oFt9WNPFC4W4ilas7vecGoX3TSh9r61oSERLWRiLYTlT
bJJf+iYw3kdhcncT+nmJ3W1MjoA3lzEP/58IkODCd9YdakdWvXbWDh2WGYTknaVHIPKuP8zxRFa/
S3LeTKwzxinoM9HNaQRPsxGHMh4z48XHaYvQwkVmy/6HSwb7SrTRn0EJeEE7F3FWmXMGuU4N6RNY
Ik1MNLfaJrZqSOwuK0QbZjOVX+zhzZ11O5nLz5WQGVsMBKSBBm7Xh+HRvARLOC9ThUTyladAz/iQ
orFHDC3bbPqipF91tpAr0vgJHYYmtmKMqc1CL952g1UyGzr4+wSPs4EUr5I+2od70DE8tzSKHo+u
8VIvMHm2rshQOh2GhwSbganeZ/5hSNN+WBUd0IcZNysmNPX1yY3Rze1pKLnjwOWIrtdqb8boYdUv
0dhppe6JhE6DlTyuPkTbE01WVhHKf67J1vuhEbfcXof6HWK84fgN9ZuTjGsCCzeEOrbe6jTp2psQ
y9BoxVlXsLDllC6ThJmDhGhT9m0nKlcOiYUwvnTdVN+XdcoCEkRUzuHZyChVEw1sQaiKCEL6b8Fk
EqjRFxT1ovvsquR+2UmrqGQK2ZWYgjw9YTadcx0ktNtSzLEKYuoH84gT/7ydFtrXfHQ3AzksGC5S
qS3SxrpTM0pWZXH/DYXCWlCGuZGZXIrSFsp0fkmqxvoq5PDC/O/Y0MEqEAoyqWda4AzheiVFMspZ
mlTXf517RTU4mxruzTgDeUiVCCL0XsDjfX0DbjJ9he0TPcsbA834g3KJzv3TjPFSLYoCR779ERkG
BPiTyCAp84mEKb8j54T6dyvs3HxEmC4yctfCL++EjmR1Zs/4T6ii10dxQNsEMfDAXlr5dgu+aQ1K
/7spejBFSWqEMXYcJSNSfHWWLlE+Urc9EFj+sEYLhQbVSWRWg9JaK2sZoAl/BZxv3lZQ/BblH3j6
svm9jeBLa7fTk1wvKyusljtjrkft98P5ISP57917oISlaZrisOhkH/viuzcnfBkpfAn0IzvOZHj4
8Du3DUpNNI0RZPdBoDhysZeUYnyRbGTPEgkJJ9/7CPOgCmK79gNewphDNmetiw89TLjm/I2JA0FO
6ZZ0ftQSyHRt+blj8sxrnBQQKbxBHrJxk/xTegUie808IO8hAODYLZXABbijDgO3gJviP0JrcQ2B
l5Sp1VlTURL237r0uKPvjMS+BK8Yu/3zeeb4MvfUsHYUAip0uKOvTG0xYIHyHiv25P+1ekl1DtmY
4JdvXlznYrzL016Vd+tO1tSfyY5cq06nGYdc33x7iyFz9eib9qBnYvuOfQjZuAaAqN9yyCyzx/0/
q4LQXihj5gvk7h2LUki6ZaMXb8BT89aYZdBXhR8yhNrhE6chTBTBwZoqhYG39DC8Q294mNVyw8Ns
Hg4iV2Oajbrg+MQc+zkIoEXAHZKlXXRFWRzgVQHK8vIYxsFTLHyfOOwSDnySVMnDGXNuZT7B3YAj
MgivcP56gllQZ3gr0dsfquedQaTmeT/DJGIbeMZXGA+yUxN+uDJfU4ixaRYiZxJosPc7k9JQoEEU
PaYmPJyhd6332+kkDubqcXRoTvR+crT3dtVtiJcTxhhFLV3r8VYfRyUHkqvD20VA5cYTfAu96+GY
FnfLVE9/grm/Vo8TtioNtiuEzYN1tw8mEWuObq/Qn+PAcGV6MBSW+qyOzvjU87q8sB4+wvT0PCm9
6BsuN9nwLKdVgciIdPTcD6u5y54DmV5KdO4+X0+HkAOpd3ZqK2OxVY6Kwb+FRtcAxGcwZG+VFoqQ
XPM+Bfgg7eRW4QEunzmaNJJmlPITVXaEM5iWCebpa5HvUuKWxM29LNN/cAaWAq3XnvAbmeAXN0sS
ihBicCl9OC0pEqutBTTt14GvrCLe74iqzyVN53mZKh2K7NtgXHZiDWrK+LitTeSY6JxvhxF3wiEg
oTwLZimoLsXTlWDt7xgUSN8pmXXPRC2lzOZr9A1njroU9rYF2dlf9td0x7r4DvdL1BkGwtZHDyRH
5iWjK/A+nZj0rjnsEyILCxpeZeIszWzc5VNRmWNIsBU9ePwUDB2G+vDEHLyW+MFQ5qkUsEYzxQZm
mZc5zmiRCiga9MwCYEIGXrKF7guTBmuIjcPLrhjcdw0BU7813AvgZ2NZjYIZgOHcPHGDFnZxLBJo
W8OguPW4H+RdZJYTK3wSgxXHWR2PM2N2kQzTgSCgYod+qaeqwY0Dw60a0PPefOMktIIbP7fmLlnv
/yNY2gbAK554WO7bxHR5fDhlsOXfFUMggaoKLnAZryjhD09KSDPZQ3YKJ5vIfAGeBlF5kM9TZoF4
s1zPdLUb5cMr6dd5cfoXT3nepqMoOOgVU3rk493KPo7T/6iruB2MajIboLmDexSkeCzI7l78ltuc
xxuh/XoeuQQ8FsORQw0rApnylOWVJc8AbqXVb5ATvexOwQ3eUc6F8Wgjk3CTuWSLgnUunQ3RHQsb
kwuCnY4DHf02TRixPC4y1C4t7Is03x0Qgt7sTfashE+pGY2TpZNS2UQdG81pgAHT2h9NbwEsMABr
EkXx6nwUeuk8tf9YNy8dtSW0QRfNxz2BaSx8sduTBvmnxR0ZF5m0gzVCi2RsXnDJYD1nOV5hF0XJ
O83gSQknRsARv4rjTmLrYix94fksGdwi2gRERlJFfBTzoE0iez6WtaIgw+07QNyluutZpmX7nvAO
mo4zBIJ4PHw3pN0DTnLc8zpyV1amuW8SClqiCIaWfsYu4M7SrFL6w7YiplC1FmUG7g6r6E6DBmdQ
XjbelJJtCXFZfWDUYk+86Pn4I8Y5BkWid3qSBF6KcngcMMgoo4SfhDpKjBIWa/4otbtbQIX9nLVm
hGGQwoNvpcP/FLHa0qSvqrppyE390NIXAtIKSLwvRXmdimh1Krn7kWQrkANKpiwWKP46bXNMAbhq
m1abNuUqhVCrCLORB9Kari/IR92g+butDWIx/VDlWrZTkGZvoxAzanuJLFzaiC+bvEEqtz0tIFN7
hVPb/S3PSZXDAIaF6+nCmplZjIl3k2l52DYlXq+tBTvcTEt6/tLfn8f2pbwR+ZYhaMXaZc5xpfx5
zoE2aX8s0SqF7YZAHtea7jRQHgxHcp1xRcB5bLsY/dMWuzXye0tbGAm6+TO2dXOUVubiodh6YRS6
W2tl5RhQo0IS0OC9UkLxndWdBhKCPy7thWvWfR7cZeWL0bh+9DvmNeNSneRfMmqxtF3MgD0EZKec
wTa7QB+I+9xfPO83AJf6Ecz5z3qH7V00nJjIWsOmMsF3Utgq/oziw3HkWNRq5I5Fd4mZf57R9sfF
fyS7A0ZhyQ18CC8BvtUzM8LAWAiNAIDoRS4izmDGPmc/qy/obwTj92ySjmOI3SxkvBvZtThVuZo5
sv3Cn+n7roMcvXoAJ9z5HoNFB6Qwl8V0cxxg3l4DGXYFc4YqcxB53hCXXYjdZDCkLOqOwzsNJVks
V5Iqs7p3xihlOvO6fRFUkiaMeMKTE6oajfXyZEm6AnB6wie8LDB3XiErhUfX4WCXPwTkBjXnPTIm
YGRNONU7H4GtLQTQsQP0Y8BLldOjSz6DuGUHConsVSDT4vnQ4Bhu17GjgEFAgJMe7LOs/OigLstN
C3Ta2UUQRMPmiqo9z0If3EoBgc0mEzQTV/AUIUDxBVFbbEyr8pKjrTF1Ejb5KRLeBvmscJx0CKU8
2Gh7pW4vxX2eLu4WsoDs86qhBhWWz7xag3rDTNr+ZERaNdPaBB9bVWvJhP8Jjh77UvJoCkOwW9K2
T0jdWtafDA1f6tiZZ6BUww8Js7s/JKrXwU8xIlJ41uVTQXbxuPtavzuYnLH6jc0DyXxsiyuTvyaC
hlxbsVDo1whYyM7m6+P2XNzyaGZxdaVMOZ6MpNhQZBmu49L6fyHebSfor7OG9uT1v9Gs1yv0i3wt
H0tMW5UvjDpgRnyaK1aveEL7u24saES8asMBWQSHv7mDJ9naMYlYAv+NqRGhEZY8IiJbfES+QmOc
ntCDJ18clL3OPoZgeytMJNtgQrHNK6HXTFYzMmbDjrf9iNu9eFOfhjD10aXKVKFs51r5Hg2hRhSK
p/zpog+Lkkwx7CtG/pf9MbgbPLcVfmqxH2Yz5XjTiGXeLgYqRPsNubjLiSiecisYAuxS/G1EhzrY
x0Gko3T6lOnj6Me4XMy8pEV2lo/a98ttnPrDIW19wL+UsHNA029nvQge76gR4w7fwlxoJQRQR/O0
YqNUgkzBQApPnhK1DCQbEGy171fQxPBZljclQGi2c0vhsBRhxgAE3M4E3w8rHq5+pxdwW7NMulTO
NwqLUWg8WwYl35wb7p0/qecliD3cSxESmBsF1UAGMosHzBLMdAb6ppnLIFrgD6cOR7NUYj+Mek4j
k3/a6PDHOpcoB9rxZgNkod/0tma7kHJNw624tKjsJgE9d0ak+UM9fVXK1dpsvaSnb6BlEF5eSwoE
u19GbuOgyj6bO+xO2GWqvOL5WCMJITFHZFhWx/tFyXxoh2XCIttojriO68BfOp7Y2H89e07v2Inr
w/hjyS9J9Bn5wIklCvEUIONRSGUecylGYN689S28jvL2t+x5pnVQMpCv7VGXDXjF8ycCeBbR3s8m
O3Tx491VAy5fFmWwah7+tWwiThvHT+6XVoevsI5V2TcFuQHI0RV16HLbBZDxoQKmdjQNm8MdYW+L
5sKWn3ailiUt1DXbu/w/Sf2u1T4MpYT7du0KMqSX2ZnTlfIOh3ym2umv8gWcEQ5LoqGKWTn87uL1
4CfYDewJPY6a5V7rcDulndofXRHVMV/GDjaFfwco39zxaTQTj8aC73HicDoCENNEL1+YLUubCazS
S9b5iYap74scnzcpiV6tYpivTPMaUz3w6+A80kAJEN/zEsKEYmHNuW3c4KQccdwg442ZJfmC4hIT
lauqaBCuImdHbZjsF6TlQmCgLAVl2rID3lJBFA7eNjAVSVpJctQchbw5UyEmwTCcNDIHaDPMmXZc
pBNCqNXaTaUW9Qtavm9nTdM0eP2qbjrsP1OsCr3uQs6BdsdCbohLc6CNrZAo0kX7A48/KYJOtFLi
vd5d4FmqrImw+gdZtef5+L/4X4uteubveIni00oUSza3p4PYbvFXimggftwjnOqj3+nrJ35HypX5
5OQM+h6xyI2tfd9RqfvSt4agsg7K2Ij283hBzuVfXAsDNJEjwZAdPdpXHycKmdNDvOzxxsPLhs4t
QCzpXJvAM1ljZewaH8i+ikzOLjJntHtddVX6e/Q2ln1krhR9pfCtuLEmJOJA3hIzUZwuWUpj9PKn
+PfPStxue/fvJSq9aSMQcGO71/hVBciCa3JkBfph7mLWPTAKI6Bn6x91FcbDX/HmUKJ30eTTeQW5
raC9bMwLYVN/NeEYIqWH/icku7n233kU24m+BreDuLo3z2KbZ2ILADtvvQNLM8yMwgmiP9IMCBFD
wapG6z6sdBmumf5OBjCDbgLCgzZe0pOce4mk1YNsCwTV6lfcus5HteighxC7PM0cUOnlHgh9Sz/5
C6i4Zs+DA5TVBJ4us3FM5zVfKB428sY92yiOqkvBy9W4cHDqUMZs6jcG38s153xN6dl4kUx3IXPX
eeTdFKMLZbsUP6zv3XeKOJFhg5tU1NqF0FPlC2tbPi/DwXMpoQoAYGmIomGF06FwdJnM+QYNLiPc
NkDEEObUEsrzQKLU5BHuGdmL5YBVR0rhougR4HBUQTgvNQ2jY4mv6AOdQE+ooata1jrzXZdt16AC
BeLs9ERWoG4WqroNdNWQgciwfWryJYQCz0LvdY8Ibl1qDGRPZmKoVLxPvuVa5urFEC8KN4JFiOH/
U9tg1q6n4yIjI7cyuoUdJrMLvtQLG/NLU22OjGtxCSssk3ktSz816bVZ/vGCbJKmVgKTu7wPDk5I
OxbUzzaMzCQXEdrilVnZVbVu9hrNKj3S4M6s4KGiT0p+k2vuMqZebV4FRVGKiTR16W6CCMsWpZpk
iw+asWV3b8FTppF4pAe8F5ji4gcYkhVAFSadEMVGXZ5hDHDKrKqveETB2OBFKRBsb3uVLWoGSxPL
0pPMgbfHYi4lJ54KnkHZ7a3I53vftE1kf5ZtLcVcUOVB8cXcwbLrwWq1NM0ej0A/jLccDJZEg+Pg
BhmbNYDXAufIFw5BIoohxVdYUx80wjtVEEV0NAZTlaI1PCV5jWl/1YJ0KONFYmeNqb+bLa13cbIw
8GTBH9kMU0Vd3jqiwz2geO1KVBB2TsA6utDD7sUZMrK0bOnNJWlckpy9B7iv82pBu2CufkHy1E6m
SlVVwo2qvXh3NGwDKAP2hT7BMm/L3RIOjXndYYKlSNF8FE2Nq585yQHGw6CbLLC+SA4vYGN+JROW
2OXTIq+PCx56KXYnx9DXpHKqLalbe9tjQ0bx36mqqFgMxnvXObESSq70mO/gn3tlQH59r7RQT9Xi
xhVBMk3QoLyEKq7thWGZaBBF8NZB7+gxd2o2hXFTsvgd7jQHKJVF0EiuC1YD3pAsG/Bf9sSoEyCS
kLQaC1VuUD+yU5n5Ip3zkdWDYefFkiWCY6wHnNAu3T76+U3/g9Zwd96ynN/rqB8mbeoctOaBzqlo
ECVy6D/s/ycx3ea40US+qQimsYM8R6s5Hdtt/qNieoJ5n/p7OaS+4mfpQAA63E292Z63EgR7w4IO
DsYPHlKHVwSpLJeGbxsrLSo+ChiHJYpyNhq7v2FtzEEvkgyoUC0baQDmcmK+6y92KeBeNbEseH/L
GVO/PcwhW8ZE/nnUBmqxzCay0SewbqjElywE9ZdVVZVcSHSefhdbhhvIXCvQdA28JRV2wqvkq3ZG
cUQcQo95DL4JlvVWnSJBo1qxF6KQhXZSqa6xUHW0vE1wdaqIE22gwqejc99zfmrvKwPLBsnjH6+y
F9/cDwYHqWzAeC5MZkqNoZ/Tbn2BPE3upMNovbW/o22EltmqxP/YyZti3lA09JyHH2CukWmfc/kK
YefZk3ZPCJWdxb5deJxhJIqzM1J6xpqrZ8cb+h0KEPNYuKp3ral2gDliLjwKLJZ54jH3y5n1l9ap
wa+zyczds+1reeVGdm65PugDch+khhJJTsJ4TCsB8YA+chkpaCW/c3Dg3M1/KNYZU9o9IyWqdNtc
VTy9DOXVt7eXuWBOer+uXNZ1aTMQtZ+cUN9lcMy4z2x40ZVYvN8E+LPv6r5eYQp7wdGpf9HJNrUK
j9/1lgmzKFB0BsHPF1bDC0HW7kySQRgBK1TY67eICznS6YomVNavhZXgvP7m0hw7xztQvlL63Rg/
luzIdpuhR/KWrg6aNNhsfuzhZHxHuGWNi+UO080YdH5PeyNKr8PnnlWGoI7YMieeMprJukXcAs9s
NGzzjMW87ZP8HwGBiRgf8jhR96PfA4NIiywum5xHg500RN9D2PF4dk4/wCd0ClrG749NoTM11Ekh
sGJlI3Voo+O10mzSyG+gnJxpFV4438fQtrW48DLf6YwIpJm84M3JfFgX7MQfWhNr1kgiRy4/Mqpm
d6WrTOVV7EDWOayiJc42UVzh51/4yKGh+iZU3NG0Vr1IutXUFK26vlNVBo2tAS4BTmTqnjlEs053
U5tte0akvvwg0bUivTcHXuycks4qo+r6R4BFiGx9ePcBWb1KDpzeR8F851cB4cb5XrWF5mAUxrOw
EpQqxO2OB7Wz5HsRcm+ExCy7YA+ucsdJg2vj64HtHApk5ayqCNCn+tDBqnDNkcG6aJxGvYzZEJ1D
PEK7pjLCPFr+I3XjOUt11dLZMOwe4vENIZ9SsbICl6LUQR9/1iTw9thJvK64vGXXAtNci/yKdvVa
IJ5zhJDITBAmBkWiAT8+6inOn9srHG9pYpjJuVaTVs8J884qJ8Iv5A43Y7WAzV7m4xl9A+vMN/FP
X9JaGWkarCuBErnhmx4+8vOSHEBdY5E+IE+TbQt4tT8AguaFF/s58Rz7YIzk/nHCRDb17wWeUvXT
6ndBUXd/Chu0WgBpHi7ib+j6bN1juQWIC9O75ALjXhcS384zEgPABr3kxdOumZxD3da6hR/K6Ay0
Y5zlaCNeTw9CTNHvyMbVkcMEBeYRmlDcVT4uGm89uSqGkrNDOoYRM8MuzFwsoW2ZQ0+SXUDdpX/3
lLonQA7GQmvJD9i/DZxfjD0dAaHlM4CFqmZ+tpfaa2+A+3BJPy+srY/m2iY95AE+JL0WoRLjdfAQ
Y9MiwG0SNbPlgNq5J0144kH3TWgb5ITnOLSIF34VcJ2o4uloDqYCPTxHPOKyuXB4vkF5itIiDCa3
ItpQkC8yF2/ZwLE01zzver5YF5T0ub+6Eq5ywrTHsb88VW7HrgO+VREWnUHrmVcmGTLq58QIGUbC
HPUXccStMTQqj9YFGBHN61NkCMD+KP1OBxy8BL3EuuAuWT+fx3gcJsdwwQGoT04qz9AeXtHtd5qZ
352wf24pgjS5GJkwgvQXH9ICYuaNq1+W4sAsO/5+uqieMSDRVtwx4+RQ2cjL+hOXJ6dv20WS44EL
EmccxWrNfpuQjnDHLtBOs9BD3TZB46C9jabA/iYqyRIQTWDvpievPBUs2Y2fyrHIq/CeM0qXy0mJ
asiXWAZP2Wo+oAqRJZ61ZBZLXvz/Gk69++RrU91LSwRqKJRGRNDEd5u002XSRzSKXDPTdB0qAl9y
gIpu9xAN/uLfxzz9Vp58nSOo1c71aaQKP3CXPF6f4rF8CHS/RzIAb3JNswWsYkJzDI5Gnbq8vnUu
FDN1nABWy7gVpVFr0hKCKRryPoDrs/jqyeR3tU6tug3t0lrad+Jrw4g+Kaa5OAUffpw3pTaw+g6X
4hmULUFQMVbbEEEzoBNLsgPwZkVSPi0su1K9CCXc6qpyR/Z02nL5dXNkrSYL1O/BUWG9j8ZAAD5k
luP25ihSyeLw2rnfFfrftQ62hSBuR2HAITSwfgU8QVhqID0VZocBoHODLihtadn4BI/dRJxr7Xmz
+9ad9LhtJxnu0lnzvWUnWoYwGqD++jKHQqLrigoG/A8tPV7PP3HD6LPNzNoxv7HPrp4AnDTmOm4u
prjN7G7JeYqPXED0fRSnM2ZQyuhcfEXbWEfxLhy6LBUCg+exZwwY3N9gs9VqI9NJ+sDd3Puiz4ee
cRFTRXZjy0QfnqbhWrUFKWVocl1RAc0bkJeBI3U5pzW9kWLMlzRk41L9nkWujOk6SHHIphvIIpxF
vgWsXsAJHAYz0ryCVBSu6aJj/EojjeYN1rusRlZKm8TZZTbsSkDKb1RLccNfUksydqJNPmvCz929
nEGALhz7xtBZjucxg07iUj9Ti6VeAAji8yVnowfVXWWq5o0cfA5HB4/+3pVJCsyuvTd4rtO4kiDN
NGaFuJUnCC8lWIg0/yDiYpPmtXB40iaMQ/yCEi56Bi+ibfDo0PM+7PoLh4oXmfiHQNLe1RAbSJkp
p0eCTc90NNHwnDtleg0UyXVQsv+Hhcs3nDBs3cJCzgneO230mJoJ5UEjkQGRsYyGO5k6SXS51Ben
CjJcmYwmZBqGbDRTJ6D95Ag43fcq27zkII55SMnHr7P/h6mhEE3wbyB+IbyvyEGEWzFLZaEgpdvn
gdTgmGskPZhY46JsfP5Mg2e916A6JWPjeYtjUvtasFZXcl0UhoJYfP8FEvYu97rnqsDFDZU/W1Mg
h4r5+NC4Mav5c1KCN9iguDn+Xmxj6GwzKIzJz0GUGjBXV6y6dfFUwOid5xSA6uevN6c3iUgPxwLK
4XVEwO9n2sFQVS4UgAvGCY4bTLdKueSez/7BaPweThtvJie6syS82NgtTF1sasAnqhMvb0VsDqRD
sgWwRBIHEkaUr36xpinuI+Fpy5onBzRMRLeO26BlRhI7nNzH1LR1JwDII6mtcrgy2SeXCN3NJDOW
r78CQNAgcy2epSnW3wYfIvAX4/Z9Mio/Lw4OP5tImkZw75nyjwsH8Cw6SodJX67kpdUalmwUpnyD
6FP/0RYfym6QUUF5Mu/6kg07wnPeqjeYOV8/vHvUNquDFUsUEIqaVMMKwdT6l2Ezg6LMt+2kUgVP
LSSb+S46bZDwWpRNsnwVyTJT6V0Xrhwuf3DhMgR7LnevAefKytd12HEK7zM6tioz1x156cbhS7UF
n1p1nKu+Q9ZJaoZ4p/4C2nffopR8LWqZo6nXNGa8/u2nDOSHw/9PrZsiHvafU2VFSu9xbRwMonea
DL1PaG2GI4Vnu9eX5gRLTYB4lD3AnYE+qhAGwmGpszU+IkOs3jvFLJAHA3RoxBO6G9zIAZtljakK
zYdLtXyPRukFBIFBGZ4pautYYSZla+a+K7M6AqPAh3xAy+/MeGrTiNBHPoc0OEvlroLgKQgqipaE
6zJVod3dQfv+S/UHXcK5Tys0GLjrjJnljn2VNfl/DyO6612qsliKl4uHq6vYnQ3iDtmGcR5AQP/3
/EegS+GzZHjRfNO0F6QwrJAMyW0I69zF+46nvKLZDxwWRQUaKI0CXtGO9Gr7CmxwyZgwnlnYNoeR
A0plE0iVidvwYqf1S6uJY0VfEiDfnoo9IFmPpBZl4Fq7y0CKRPSaXSszgFr/sX6jZFruJ5ItWr56
9Lgp8kTBe9wwZHlTFIna8cLsZNvEoG7gP+4p2ayG1yHsvHkk2BbFXW4zaQbTsaB90YGKWEJBxIN3
YOvqsqz5peNTQx194X53fG+re9Gi8qajVoy+xn94SyKdgkRrOrnXdIUBkRwbM3Mm/mUzFNtfuCA1
TlI/Lf7jVbuUkXul19sWHKS4mf7XG0uEHnjc80qw3jrKBevggYYcXsVnwelvvYjgm9XIRcXXj76w
OUEy/dZAC53ro8w1eTSTUnAcgrdbvbZF2hvVRHcHXmpRsyfAr4390VghoZQDiWALK/Ezmjve7Dc/
A4geRtlL+LKB6aka5d+Yv2mOgVMn1PRqlrkcgjBareFQk9Qttg57KXws85cEgHINHAnbsMcRMBPK
bKsD6/DP+pN22U5MNmX3yz37EmAAg2xYkuY7VVqnGu6VjLfk8/FKcKkJ8lLe0l+8aLhNMF/XqXAA
jzD+Tszdzdvs6CXEVKBiSbnwnIz8gjp+8jFQeVJ3iX5Asi3SOukNq9eS6jmEDDyiToQDqxfRaiv1
DAEgL4AobEAQ3s9i/z5472D06UJq+N4eYo+aPaECclZuUDEOPKeZ2ntpecXwwEqrE1wqTFpkLHV5
jTCaQURbXWJzlIDw89vAe3yOGQoQYyLpvVd0q8dDyNqJGgjsKQ9z6yylCivKfpBnzGWTFa0qGjlc
14/xQO5Szf+Da5khKdF+gkSbuc92K9lzGIBUphvcpp1bdpbOnjyiRrCZoKtZZdqSqumSPbOWobge
b+wu36tWSksMXFVnoUp3MwFyeFEkaw70bFm3YdWnqD5X3lVAuLR4U0Szdkw0WJvoG+OZAQqGLGlo
AAxsCFyztrDlxCILy+CoS2b9euMXaJqXC7lqh3TVmAEidsirCmCa15MbQqrXvnWYahSktQdxaQmU
CzHAHodiNrdZntgIQzzNCNbvwQVC5dzsl/2SjbwkN5JhfTTqyQ7fdXnKv5XRn7PSjAIoHGI1V4+U
GcPw554Cdp/6x7AwcU5su/tJZLfvsjiedryVzrYVj8QzeT44io8ZAxwHxX7MHkTSS7gfohVohqUH
piUpiVAWmaY8DK4ZFFwjhUr/ZIEIVoZAcRMjkqpzcNuLWcH2jMagF7Pz5e78G8INV8wHpH7REOKe
5cB7RPw35vDyXWZ5lixH0eOFfLWCONDC1JSV3c6HtjyU9JUkApFkgLW+8O9JEdJJ2jvli1T9+Kxn
TebJB/DiL8U0L8SU1eWQF+Up9VW4yv6su5Yr8t9hZd28KTv2DVAdTTgiwlqYCTXbzNmYSfNms+9m
yYNpRJTXDAy51nIcgjm0ykkTZF6hE0Gx7+PPZiMeW887ayvNNWY1zzsbuOJvbQVP8t3jRsglWIav
iuFaHuKINuxKB3Totidiqmd4XY6Tv2qAt+Rtko0WC9ns9dp4ocze8aLSSWtj1q/q0DBl9SGs0Q68
J9DfvtfXtj41V9oXwUhf004L+khCrLIRaF+fmSlGNbySvUdHN5itnhYioYHQOd2aq2xQ08Ux/6Qy
6bx2ATrAU86rI2GlV06BHewNzMwDAzn2UvXv6TjMjY2mK7zhq+2Lp2UxcW3kmdq1iaWD3JmNPlWS
yt8ECFnwcBxmPiwIUanmT4jRM11U60rB/zcRypxh55WBxlgzNFnYi2GVVSxvp0l5jEzWCoya+jz5
QAQwn0GPFI8sFVwn2cuDVEPG2hfeX6tNHeRNgsHSEr0z/fVhbF7Gj80PejYJLEGZ9EqF6E+52oez
jZcb0INzYkXKeZmaHjrC7W1Q1NfrSgQxOw9XECxAXBqZl7GeVN7Yf/H1hG3V0Of/cdIJvNP1yep6
Tc7ZcWtmLa4ltpdFnTFutCBJUtamsrcCdTmamP1OJZuZI3kzNIhyVmdyr2D5OiLXzD/+X6Dp8Uqs
W4mii0LvSiAuiHFIxZ2wPZrjJbKjvxlyO4TJ2uPyZbVzo1nNz0LbToWTkIOyF0JtCPf8ppMEC48a
eVQedsPgJIKy3nve4C6lzj+lDL61OGSiy4qVE4MmQT4WgZwbJ8VeoXVT20eomYTXV26v4eIxDByl
ZbKwv/MpILXQF2W+1ExT078V8ASGH9nyhbtz9Ldwcnqn0BQLhe1cBo+aIxG3II2VdsvVvHjI+XAR
svG1vWpcCBfSQAaGx44rTZ9Z+Cvdk/N13RHc+AfrVmW+/0s38P4MrxUObf9kyzPvse73m3zYeSZb
4G59nS4v0m710eMOLTU+kn8KHPl+PjOfpGrb/yo5IPAAzIWmQS3E7vznYPJI24qYDVG36gmh1IWU
5F1O2osdWBzVHsvd0M4mQuXwkEtP5pTzicU6DjlRsmMRFiLp3YkGOI0d24tDUOM6qSiIAYxdKoX/
h6sLGLQO+xB6PGz6PZh9HOv0KC4YQSbVrrpiENYK911x4r5/9UKNDVdCEvfZvXfuRnr2txbzpph4
vYNhdPn4F2i53pPLnRrWV85s4VOLmsWp1wuMNsiVt0O2Vu6biM5Elny/vcQXAbNHp7tqCfyq0+qK
W2iTrAwiQpaBgrdL6IZjL1ksql0RyroWIX6cepfaQ+tZm/LO0dKjOK6NxPwTXo1402tQoqlDEdwj
9KG91qD4dc3ou/5U9QblfXPxd2c8Lp+NnCT1P4K8Gy5Q3pP2mL588So0NP4l0US6Kw4J9URdANgQ
2l2/Vg+RPwLyozTJ1as8q2xBHXEk0x03iaT/RGNH33+sqDtTgk1Yr5fKNp+vB2hqAABGrB1Gzdjj
i3tCYD5WAz3yykD8xDqOdKG107gBfIEsl2nKFSpO3blYfgW9p53UslKdcmVjPaElmv6dl07vVY4g
Gd49eGNQuaoW0M4CEaErm0cAM6yAW+jXSpeAp1Z/Tm2Tp7MtaO25TaJ60L6Ie6TJ4yxb8RS61dS9
ES9PMPe2fl/ABtcHQ32Q1T4CO0VMm3CWneyPfs44ebLcsMo0kpyoGQqQvw+6xeflT5ghXWAEAp1K
3mtdPMTFbQ2zG4i++QZci45uZ+iaAOru3DY06Fs22ZT5vVsYOghWvclyCQ9VhrMgOq+Je780fX4s
ynQmsCiPexCmjz6sbWsVsRWpkrPgMn+ETtmDKvv6e23Gazt029Y043pLPWXXo3j3TUboU4Fzxg6J
r4RNp9t3YIC3H2f7htI7iiMsufUCW+cQYlz1igkPEW5gcOQJ8tWZYlRzNfnAuDLzrVVxxh7Mz8v9
eeJuFdaaMh9vx7tDr5weqIbe3Jhiyzv3nwJrj3jkE3s/k71rqgTMcxM+gTqsdC55lMibArxsyffz
SX+ta0tW5Ax1fv60UXpuzx+J+q6UTWHdwJliAi+gC9Q9CKi16ajJ2kAFcxCEeGiYqXU0yKReGcxE
aLVcSCMUmGO7XculenoGoYI66PbInJPS3Uv277N7jCy3tS1UWzsWHxV0TajooYMrNJC9C7Su4DSb
xhmGNnAwBXU54ZkYcOJrsYsMIkfblHs1OCPhaiLhz16JJrkn9YRgkTWlkChLSotvzO0WUN3zHr0u
SY/oUh+NSrgQY1UF9kkvI0tKtwfStsJxjKP7BcRRo9CGSEU7p4U8ovQGNNTf0ZMxNSTmX7Y07/Q5
EGL6BKFTbZhZcWio8v1RwG8kE/Yhm7kTB4lrNe7gxfJ3UzMcWhLI5Z9ETA7XMMlnPrD7yO0vByJC
npEatljqsXOgXjWrLXJ9t7rYVOXBfcw1cJO9BjDDpCgbXTBE8TkRTLAyZMGzrl4ymqMA3HEDe7sa
OY9aFVXjO6G6/w13trOBN8MGpIMaSRUOxKWw/5m0olTQkPUTn3yMft9RLzhmEZErUdDt/wa6oaaX
dR5HYnHOSmKAAS0dS76zigPbeELx0bwccUsIISKyfPtl7kGdp4epkauPrQ7Y1B9lfvphDgxuWoHy
tBDQMoaVPXMUujjJ6Ll9sFTmqsIEZR4p/4HZMiyDo7eZJF3SBQt/cMb7542O1EzjhMm+BRBD+IZk
R4RGjE1nfK8DvNEpd6T4DvRVAJ45pJtFs7K6gmDOu8wvzwtr0d//ptK70OjuWB3d06c8qbIYSUDd
Prp8VPAA7ORMNDYaFl6zfP5iFJNFTDor/iLn6WAryWbK7UntzZL5cB+EKw/ZUJW4HmM2jKKKspQS
gnLW0wqOcZwJZ3gu6UPnrBNr1tBnkWTafbOHNLzKnka/kDm3AXq86WU6yNqjK4TH0Wq0dRYdHK4Q
2eM3BgXO95lzo4VtFsmWLvR4xXhSYmZAgdJokR/mr34/K2k6M7ZnBz7iIldpa0hRmhkrWqJdfqLa
7Ta2lAbEKATYxuTpyfNdwfj1E8U+Ws48McYn5gcSFzL3O21IPARCALFbrZcF4WuQQgmPADPgaV52
qdot1MYLOjLJb61qelxL7UCoEIIzMa+ViCya/JI3CLr356fpfuL088LjvFn4BwUpudA4qEPRnH/U
dI6u3lZZy+fdGZRiihuWqFY7KsvF+wu7J4RFGk8NFz7bQmitJDNVrFmkMh5+PlasJffNZEH5geA1
ax2AMFJmyHchxllkahkUEY0ll33OfwOvCRp5eDLjlr0uAzJZVE+zz/O3xDbjqqi27Y1OyuPUJj1P
SWlYB+1aV0lghZVMrR+ienyK1FPkbvVdzWyikUdMQ0ZqeND4+wH8zAHsb9asrL50C+zIUeEjXHQH
WLVEU9rki9j+WFcpTF4SJWsACq2LISxMsG5iMZXG7FDIEUjMLcI8wjlRsBC+ynBY4sk/ssm/pR3g
V6IlG/sVyXJ+fBUeNbsK4njNlYKrg0+bs6XqTzGYYRyACmlN10kXc1cv2W1GMKfVTogd5GPKHgzn
+XdBVe957RX2iFE4PCfnxxV6qup0L3Eghl8wwtbJ703pq64/kXwsP1QVAJnOw/Gl7Pa2PR526F5H
sl+CNL7jGoZGg8EIV76yrAyiNxPD5KFoWBJNzF+S/4b1wll/qAizlaiNy0yyEAaMMgQ+GG69ZUHe
hXPXWe3w81t9a8PO3uYJdt5fD8tqZhO93Lu8medKUjp2Sv4f/JDGU4TSKXIs/66FNbkq+nTqKkyy
mEm+lGUsrfja7I+kSjXn9x2aCoveegvvqQYaTf3tIDAKzjQt6BcvOZiQrrQXyWomgyv036VJFumy
oml6CASA3W+nsr2Zi4KkLK1RYx2KI56VhpxfpLzbhsTehNyumuYJEFPjrgqrdB9GdeAIQCpqTWy5
vxWQegKuKYCCsKVZ0YiQLRt5wHG/q8PueLe0WiqGzlPRqy9Yd/ehzNw5MhDLnGKmlFLzMGGF4byj
m32X3NVQqZOb+ai8DHLbDbSqvrCZgOUyRsvtHFMItJORGJnwHvgS9/w11smq/3z8iw0y+rNdgJQf
xwiKPeFZgvM18TcnkEns/6R9HQ26wyS11s4X4dq96d1XVuckfxxmMw18GP4yw+qHYyUN7GQFph1r
+hRaae6FuxcaYYYUm6fFi74ovpCgC5OoEPXR3JtjZ6vJRnilxUC95YCFMeeGIu8Ffcvxh7Q/Xa48
uVQQLpehhUKq1e9TyuoHCYTWGzVwCpUK9qLJs7fIBEtVLuwYeNP/qXm+2HglY3WO/hIhoB+L1sfB
YABzSRs5fnVHZZ6ScRgkba4/4lEsWbqhR5J25Keyx+2Fp1qn+3rpUqGPzaFK8J5ttzBnBuSQWyfT
gOrFNYFmucurpqJ2sdwQIqpRX1j4t/XBhRZzClfNrqmBS6PtJBexvzsaruyD89qQU+8q+t8r3luA
va8e5jTrS5szSk+L29SEV1mwF1Bmg6O0iRamNfCcngECfvTLP7pmiqx4JBUJa6j39zRW+drCoJ13
ssaYSFCxNF/EClms3m4J3lJNAewnVnWBxZb1MOLLa2IWPyjmEHLpSoCUYMqD7g1l6+vzDN60+bYp
7Zy0TsEo2JSiVxl8Q+PaxsUupT/apXv1VA3rEVNsJOlL+I06QJet7Xof7b9RuAB9SAuiVsdZcUB7
AtjloA3ODv3IPVu7Czjj1S6+TSA1ajzf2t7VKo1QQ+G47tW8OLVfFV2/pSS+echEWYCpOCiEnH8C
rg3WL2ZPaMQMbSFunUO2M3dZw8LDrqfM2hDpKph7psFfWJwTjKPxQGsfjusQHZmBAFMxNmE866t+
Fch/8R69kw18egntZnv8e5ThH1QvHQXZGkjFKGQ8kWQmcVjPAuhwbSLsToF5yfpO0Mn7kYEnBPGW
LRyGPVg/4ZX5SPd92zGkkJp0LN9ZJk1+aU+nE8Ld3Sumu9KIU3qTF1GfSnrwxH4mtdfuxs821KF+
A8bSf+V1Y4jeCPVlCW1nSyH+kykdtSTTpx7zGK+aLywU5NigJ5fxj9C/ITkKIvJrR6Ib6hB8MGs2
VozBWSn2ieUxwOt3OD9AofjxNjJUEgOIlnzcwyGpF5laYnAlbwQrarjRtBd7gkP3qvU7zC9CZYcE
WeMm3slg918Dt4yp3dc6mcXazeqnYaBM1MblLmTT4uVlo7gDc13AsPKLYaiP/55LQ/ZJxKd+RxCs
N0EyX7leFesOLKC66p3JlKwvwQyDrTKlr6DpRGCX2TuKHEk2sEkKw/u5LcwFu8uLxnMM4c88fCWs
e1A/eRKNYxziNlE3X13KCwO6f1rD4kxHDyYQJak54s02XXj2Yzt4qAQTNxmv0EKjgmXIwQKqCMA7
sfFmQAWWwgFdifs0pdJxsHh8rvcmWD0L5lUqZuexGSPlMCcBAnlGwYCdSaEEeQCdECH5IOFrnIpK
Eh0LHUtfMer8GDhSi9xr+vVhBmAJywWuJQr1hRu2BN+I83GSQS0Tt0K1qcPTi0aQ/wC6bnNGWLKH
to5/UnQuliZhmHKzw4hONa3pLUF4M6VKRZ53uBy4ANnZKNO+V2XFR74D05rCLTTa6p8fOkTS5E2r
OpDxWqjt6Vnw/P2paNzrmfc8DiWW6OYsxhh6N9IOPtNwKsRirU7ZIt211UQbtFf4nGtjXAvO7z1Q
efQtZcLjIT7qn9BG3lx2e+EUuwR8ovHuIBXA4/R7fM37Vbw8juDfWWAk6hN/bQteDItpNrNv2sI/
AQchMkTSFbxnhaizUS2Y7lX5Aw7orLKcdSNPLtX5f5hCdla5VmO+qVBZIvcSAtymItpzeJIzSJYK
WLQf715NJY/wJyGxKFP0Q0geQMdq2/dnHYba+C3fwVbMirwLX0DdVyZiGily3pZdsuHy1cJh1280
7JalfiUa/npflMPd4ELJYMQHVzeIQV/x2Zdf+MwmmSiiCSmjPTrlXaK7pNr6tNQJDK1OTXso6uSF
Pp367jfodG87izFQQ2QattOUjXxkmK48AmZcUgAlqjMesA+Zn4zYIOpPEAZcDgsm9fSk3iDauocS
20+2ED2Sllk4krtqNxpxoYpPGVJe8mh/ojEPC1CaDlW9Jh0guNFONPpReG8GUbmY0lVEunxwpwk3
QyMpw5vxkAzuF5SZEruCYWwjmB7+hwZRc53PnSgkK6dgJoG5Gpe6M42wfphQ50Cgk9ECTseZZd1n
JghxWtw7tEbOTpmXe0C5vOB/R87A5+1Md1l+wllf8LLKOCeLJ0gN8qjn4qENVe33QJzHhOnhehhU
WnMS04GogFFzy1aXPFg5seLKPkz+LquefnmCS5lRl4FFrFNB/F2Rqn4BQxbep/x2AskCeI7uAri7
HC5LW4aKIf1tTxBqI+xuDPs8Cj+5mILQz9Cd2IvbHjHfLXqUK2P5QrjnyP8Rq1pkGtVKdAaLAv5R
d2cglouzEIjTNR2itORhceMHdowuQi6jsHPgSQJMiBH81X6E+Odbro8DEJmkkoaCAkbDJjDTQWl4
UfRIs0vIfEbTxm7ViNu8evXR9/q0GI4Z07yCX/4PZxcgj2QweMZEvnMDo2U58dO3b7Fwghj+Qx/B
0ClAzJpxcMTEnnlZVDCqTY9A5P2olCU3zBLhIiHhI71MejN56963PpxwyEaac+wsXD53Ovzyxu6f
LmQovsSTrjMl24utW5QR3GDguj7glKinff0NlPzl0qFHVf0Yp6hOPq6eSnUZ3rxF+Xbq7Hh8vyPg
MiQ4N9yrElLWmzdz+R3S3bQOZYADmPBRV8MeONdb9UFRvUerbAUP/ZaTd1aPHYl+qkKWwDGj48w2
rtOnJB61K63iEUs0+DoagZslSkgRsgNWDaXFi1KnlnixPphwnE/Yh59jBZER+HOD5mC4CY76fDJj
kAG6XirRYr7rAkZAEiVb+x7DprdNGKH1yRRCXb5vYcCpR7uY3yhq/hs7smCSKaNMGp2ldVH4+W0a
zYWGvBP1g0s4tm4F/CGrqatahVN0uQuIBnVphGOmPWrDkvN/FX8CbyPicbYD/PPTxljTkqcRIx6A
wqzUQ6G8NK/JU91zoQ1Sgo14Q+IpU46Fl/b6L7ZlQpTLYGezNG7F93HfW1jdn8l1vOiaJwjj1fD/
XduEaw+/+mYmNLkofwhRiKLhxK0EBSMm2jZJy7e0Hm+8I1wK0JAhIhQF5L1w3XHWfSglYQ/b7IDt
XhHFmTjezt+pC12Zz2fqS18FKl7MyzXnAf8lcoTkyC2guFghqrJqJ7GhOTzbImQ12I+7lZuqMS1b
SUSKC3G3+BrZDXvNkwm1aDqrSy/rWrb2Nuek5hhNu0ZiqHPUC+0HL67C2ZIPcAVFStPTFx6kYZqU
/i3HiVY1qTatrrkRNMo7es7b56nqoSPj1HGvIxl7+acYxKNdPMIUaEgrY4ywVc9XrfR9n3qrq1R4
W7fCw13ZQPweo5Kn662IYbPk4J7QNfbAU7lqRe0G8IFkwsCm5ehgPXJn9XUpEWY0l8egObwCGeOi
V3i8nm9niJvTuSz1c+pQ8vHbJblDRthxnsNjDDvLx+kWyg1TjJ/QbQbp8KeWp+ZCDT03VhsWl/OT
XiaNxQXXk6ajC8LeTdZaXpCY3hCfIqvdOFWpP+L0e4w7vVYZyk6Egpc557AHGgVH1g5hP0CTwhzM
P0Q0lmQy5C20wC67XxKmzUtNL6ytkBLeQJtHlB73IT8WCY7T3QcTY1OXDVG/U3j2ObavAr3vyVvM
saRjPLYwNdGyIS6BjjjquyUFSwqh4WbqkmQDIFnnNpkny7f41vKUxzpFIV+utMJ1fWndIxx/DCX3
POiPNZ34c0SuJcosZXz7+lGbZ9/PFfPuSew3VEjTqFG87qhb59lB0F6bmKe3++yHtO0LqEgXn+F2
mtr/yfM9lGtNr6NodNR+S3ihbQgkGfOADz5P1b/RvQhdxbSk8RyRY2BbFK592yNK87LoEF+0ozeO
bMFajqfQQj8wMBwi3F1Zqpa5AmS8wJ/yIx0DBIf5ankDHCCj3pvcnEZBTqKLcotyzfpDh7byI1ib
lKOscIMZLRO4oBU9+/mPnLM4LmvPMrZSK1yzdpvcY4SbDZyLbGjG06csz0HVr7VrlI1ylBPnMKZw
Seu7xaLRS5S/+7U5JU283MGATxdIN2G0e/XC+N0NupqsCwSU6gEVdSweU54Wz+JXSH1Tc6ptNWjg
k40mFYtY5l0p+FSGKVEhDMduD1zXj11dRAZ7Bm9ZXmNP8/LSlXEAQ86m/xaJBGdPC9cIJC6ItoY7
K+PwkuyrsUcP0W13c8/lrLA6mEjWmlUHM7qBlE86x9lybxnAVEY6UzPUtiWvVRfqieB4GMCsVp3L
QnM5q/6l2DFZzqj+WXnVHiEo/D8WuTuIpsbMtgZZvuxrYmfknYdBWFEP3k4Dc77QEdD9qcDwfUi/
PMlfOBSjHBSYLdtVdr8OdTWobmPqJlqI2KfwpHxY665ojfPbgx5qazini+KbuD6n8d+BYMytJDIP
bzbPX9uY4HGESt332mzixk4dYB+GIigaryodY/gYVCx7eljgq9/zuHo6nhxbQHUG8HlaglXee1S8
JdEOeRgeKfXmob3p5fBic9WQrrKavfmAZFqlGxI2hNrRWJMgfRv1xyyG5kW10gxVXjErhO7KvzUs
R/+KNzRMizIOtHpOLd8bUF8B7lZ6JqiSJZiEI5tudaLo+iVnbvWL6vOgfbP+T0hojeIz0c1nk1nZ
p5JpcFvhSYrAVi32cvas3lw5jzlkOpV49qt+dKO/i3CFFxcDpPSMq2qsus0DMHN3Ly3aUWzeyURs
xBhuL0iQ+A7qtAkj/KU+YkGtp7NTEN3FianJcetPqFV5ZBE+b1JP/Je8mKRI/uNyy6c5yfLr+xUg
CPhIRdgfwpH7py11j2B26Wa4ZaX7cEOe4LgT6nlxWbcqbKQnWKKYPKXI0Aq2ZZHoiixpvB8HgLyB
2unw45AkfGOBUsGzb3pObYr5wxW4HjwLa5G6CDhUQaXJtWH+9EWq7r4g61RV8Acb+GgSvCHNsAqZ
X+UmpkCLdzj8UUhyq1ePRFYn6pEM/osqKniTsGwCyGn28bjmFCE7M1CtYp7D9PYtVtf6rxOdYa+w
JSb4DkhFE1YJB6nrfVXm4aHecWAFXMcqOW599ofB/W+lbO/jAfOMjG9LjTR3AIKsl7j6znpdBTZD
QDYVlYaCDgArsXIK+dNuAmWU2ZeB/dm4qCipD9H28wIMhSaq0/ssQD8BpmcLFNWhDOi1uVP8IlxW
tQRh3niV7OjfYTw51qqZM8ARkqvgP8A3ZeHm5cxvdflbG7d4oxIHg+omPV4rr2aTRQ2m2vRsv1TW
c8UQDF82AOWF+2pAVbSv1tS3xTW0gW8P8iTdTuMrQn+iL6LxWffnf5K0lXchk44QGKdQs/DXn+o5
RxEfod8il7m84KtsHcCl6BNbmCiL0hUAlF4rO2UH+l++gifPxvnr+jZKJp0QyzIzA42Ij6541gmM
OfCHFb+sZ6JUt/Pz6T/NxT1fpZ2En+QnjwvJRZ9z03Sq5HuV+gRVy3clplQhJW4Prp/O/cUAK638
bVlthh8AUfwG/YaThvikQkYBD/cOKpYIhnQS2yiYHQ2DwfU9k4GX6/yQXYOYbgeF/pjBg3lypZx2
frt1p1tFgPchO9Y0j9kbZUUePxozCMTYDFXqpoLrHA8LNd2soY3l4+xpfQ+DaaVUGzCcbz3YON66
mlK5KPLctvuz5J5lJoW1JwPC+SzGntOcoAVHEhnVEBxAqLsvIUfO7Yz4kUAnI5ExWLj5ccLpHLDA
sItUgb2KSuZmkr/ZHucCqAL+Z1iYusMucW2+eMbOubMpACXm6f7QAEz6FB3Zp0QT9rQFFvcTJznb
Ufp76VgERZLRGScJf6deb/wossWMGm+z6c1X5BJjB/i+cJcRpEr2GISS/ke2ML04yFLIEHvessbl
Evwtjs37qH0goJ3B2aYqidaa0Fvpmas9X3IrxmP5YTZG7gu+tVfDGTb0AJPdUMn3XCmjymxIAxx5
vBq9Bi63gQ7Wq6WSX33t7N7ZKUUN5X+ikkLKHfp/xTMFbU4I/iUZfbTw/w2SrTZBYpwqas8wgkbq
7/IKpD7G0zRZnswArz4PwsOpEIAqDB6DVpR6HMvv/mWMTFyIQsiHK9VsZ9PNay0L0X5y5uU2bq6Q
0N5Wyjl5qE8SR7he32CDjGJXf3bjh9NLUd1uKh5TemU6kDxBpGl+Jar4ZA+HYT9/lx/32d70UCGg
H1Md6O1FYmRNNZXkm2fS/WH/i4xfzWxPTYsv7+9yzktwzdbvfvRhtF3WG4lXQ3y7OXe95bBY3txs
IwYN4TZ4V9cI2ROtZMeEXwM9UP2AcX9WYJlHwfUbG76eUU59PBnxh70QJmzmZVvaWTPUfVsD1uwV
eWt4t5ZDigMLGYotiUaA5lZDPr0Azn95GJO/IZWSaJBX+cZU8gdOV/YA2aAFa0Md8Z/+ywKczRBS
v0dqVJ+p7zvRpMRZbtub3J/ZMJTe3S/xTOZGNPtSMtMXCZSblD3I9kpFVLk15SGcp9OCDXJKXvkE
J4Z8kReXeb7eAGi84QZm7Ia0Np/3vdU7Pv03nuEpHckUw0i+PhjlGDwy3AyvRIZ7gQo6YckqEMu2
uCtsjg21sd/iy+8oFUqFn41q+6vxMHlb1Rhzcs3jnQHmj7IY0G35q5tPJ0Y+jQXcjZDKRwuEb46C
s+dPojaiRyd+qLXW8MaAJokcLBTZ8NT4RI2hARPoHWjCGKgKMEg+GANwcatRKh6ttqGw0f1iuHIT
M4EqTWeiN/q354jCYGHnwcCuytUOTsO+svPY7XuK/eBzQ6ugorCPIv6VeDF0BqcJ6yEFFpm2yBbs
6B/2iRYU7csy9SltALruSi6bkBzvqkd0btZrvfZBOEYoKLg/bcPQy+nG9VRTuMD0f6SZKi6TYcRg
/0eXAf8PCtxv85QoLyANQimLYCPOTwNJxoJPol+p6hL2NHyKXrtzxEIiAWXin4XgyldcXiqqca1W
Gn8JVXeQw5Fld5eSn9d2TalZOgBmcdw7KUtg40Db26yBjN+7VnQJTBUCCHrxstL3/kPsv/81oIJ0
aMnv/iLLBRKEUKme534FLBBmfkm9oQE4+ckLHis2ms+i6oAedRaUqX0wRPIUtLRSexEDbV5PrxtQ
vlVTRgSsO3/zxG0IjDwvkGbOjw2G/Mp4fuh5zFvnUC4j1g4U1RmFcGxaU1uJqtA8uyn0OCNwCBFw
bArTK4W72foEeeg+3L762UyIxIbgFimSPyzTG8c2EnRSJ5Z38srzWUCabKlKYXiC+iBWUmjWGYL2
/bhrN8MPjMmDjEKMu3fNxilW92eTr6vl+KFnc2FDEq4asQlti0K3IvdI2zSEB3xV9nWaMNXmti6+
io2enoNX/iDR1p2ARyiGlqfV9hLjZylQxjSUWaQY3IxOPERx8TW/PlW62r4wrF9rig4SV1lppuWb
oUzqMHGJkGJx+n1Vlq3iqnC7dOz0o0Vt8EkaP3nHsonL+Kq/dLf1gMJQa3esrepu8yq4byxZmsfZ
PaNCPpC6l2cS1LzWbg3P/MC4fyfrlcZyih5Q7aL0y9Cvrt/6hYmphlzQvI7xfUiuJHyirTcEQuPa
RdukV/qmR17YFUNZIe/PjtrZIv7JQtv6hDrt9g5eXXfoiIAB04Wh4wfJV2F87IQVGZU71sa3smM7
GEZLz8p3Deg7mgpv77GqFVmBxL4GKphw/oIOVPHzCrWOB7nswEeUJG0ZPsjc6UdWRLpAOFo4uDbz
kPppg/R2jIaM5Cng2VijU6YdU7xSJYcGGcWI9TO7tLDfROxxb4egxUirLC6c2I76/iCEj9E+/fTP
/bMvqP3myJZX/eU1UtibBG2aIpHBcmFM4jkrjcU9eBDuwGXdgxww1ymLAXZxe3tl7WmmI0Po3hdo
KOOFE1nIQSy7i+UqM2ipBI7N+MDaR3Wn8Z0lsE9eE0/Uo6I2bPcQ9JCL8H2VyWPQDHF7loDcwCJx
N+8rScNQh6G7SoL4JhccKmea8DABBE/9OdI6LaeSoffbRc2gJxuyIF+/S3wyPxtn/x+wuzxyCSeU
HxbRjQ6Ftphq4al70HEdfbmebW+RQR7dUacrLUWIrBLSNy0ngTkrgLVg/FPdrPJ+8X/EfBem7BcH
IogCByKVUJUt8nw8+UpmqmUr6H4e5tw89o0SYQXIOXNDlc19pTY9v3IRbOYqomTDmNtt4Md9OVbV
/tXTxUB3Hg+HnNW6/6bwKcMSFV3wZXwHD0O51FXfRMLWMHo49q/FcrVjTmS/8o08mPA92WdZqZK3
WyI/gUncg2DPWhuNnwYei3YuEt5AZWJ94N8x8jYAznos/Ij1Nhlow3RAiYyb/feiRadsewBWTIWE
f9yqw92ablyAepLKTbOlS+ZIj2s0weQwla0wdghl6lzZdHFD8k+zrFdHI2T2jDfsbMTdRz+vekhb
fuSmCz6vgs/rsWp1rYIenuj6UasMp7gd4jiql6JdkyOT1d3d+pjhpE6CBJ9tEWLWD+8NmGtvoVI0
oDuzU1sry72RB2ypGitiTESErlQ+KpF4x74zSn53U+XhttiHPWhcV/LVJESG02ztNXcntIjVLbR8
QMKViLosdKIlFO4w9oBgCj7VhiGWLbCLPZorRcmZGxKt6D7xZAHF+mlydL260v2clUurqAqHpSVs
0bNTImiTiK+JyjUIdRxVlUryouubSnmC7vS6k2s9NcrOacn8A6WHVDO8zafcSPZF0dxsYLQXu/ec
CLtcqaJ9CiESmBu6jG6ncUNOSoZgMaT2X9jUis8O7bASXGAFHlILeeZR58P1ZRdU+DBANQ0zTNvF
5hOT2+nFuwZvLKaSjOIqk7SCTaxw7oZ6OQXaHGDZTZ3Nl/C9Y79cAJR7ITADI8R0fs4Cf/Ip+eX3
/7dqbsn8r7PasMuQqTbb3dnwx9iIuzKJEn1nv3TOD2+hO4oWrt0l21F6bvyWLCf330ru/ttqoC4d
0VOY08gv+FVWpFjJ7FJgPwG1xhyQqCNZKtDPNvmE26mxateKqlrP7h7ytHECW0E/F435Z5WBGgO2
gZihIVWhgaCEkJIDKN3JRxxzbivZzzkTaeWRSFvPyYKuC0L9RtMUxQyrvigt8K0g7CcksUklmqEw
MTYMTJiPhQgD3RmKiMrvLRiiYVhntTFe9iSJUe28L13JojUVTp/SZtmCJoUE9ciJmEQjoDWp0PsB
CDV1/CszbkqwxzW0ylaFXCfRBUX3ZORM41wwhVsm+iQUciEu/O9Rc/3ELmexUuNpVFOj0DkRAG6u
aYpozIcDE9zLHpYd4d4HrNG8DDW7K1QY9UgnIp1DBw8wJ+VkRGEQup8udQ5KXqXNhIz13ouVc9sz
9jq55Ou6dQGCyzXk7HPq2s0cViFaBQO0+Rr8NaZ+0QtK/x7iOAh999oyVzVHzj8lQwhhQNdR+mZv
PQ7YKbrsfHSgS0+vKvZ3lGctmwKxcTBy+gF7VseOC1xr244XoaYiWTRXcKZSY9Fz+ToJTGYNUiNM
7J5ystxg4SwbF/x4eE8TA0FjdTO1KF9qVOXJSAHXwypKbWIroq3CPuEHu4hTOi15c+9v5yQm/Dq8
5wcpo45bJrcbw1k3OKxqIIMwSXxDowkh41uytly6CZ+26FdPJE8sceM2NYBwG8HVGV+d0WXsIZta
hjKOSP7N6JJjKbs5o257TUeTpQW9xUo5da15ITw8HnihQsZ7oYd3kSvoygHpQ4qJ7aYs1w/2Ozre
HBKfR7Y/k0FjQnxvqWrIFaVZaNkYYl9Kw7kEdHK7xBdz3lmmUqDQcu6ebJeBUjs13cad49HEL6C5
2ojeLUVgtASS6t74FrRYJZMD6KfN1Uwp89pZ+QFHZA/uQ+bndwt7XiH30VOrP80fu5u5/NVEyHyc
iTw2ZyYgqMmW9Jmxab1rv8KqbcuACLjPaDZrKgOEFkAwEPmbdrRPKnRkdquGE3K5pH1noCfE3fh7
7sH+l3odnM78iIihjikYIJOV1wi+D7ySpBNSGCXSnyJNxeCA3NpQmY5Ap/8nMTuTAbZV4PEpK36K
3kt9aoQt/cNBHNHj35hw2RMXKc5ckhI3FPeOFVP/4LmA4xsYVVOgTiP076IiBALvftc7ujbpxyBG
ivT/fwqn4jG6zQg/M9cIEJ4g+Ln7Fntt9Xt0547CzKh/I4gWGdh3xPd39xwJSbu0a9458NVYSohh
yzlnHbsLiQ1U8+TilVCE4fsN/3pMO9f9dN8T8ZjYAsc4llI2W4MVH393SKwkyRobYkyp0mGMFqg7
wODeJGFeyDYhAzmYdA7WUmBQ3IXLxCvUu16LNQCaJBcICNbtwxb5rD4zD6ezpOdRVN7CxSiN3B2n
4/t/QKlqCleJYpowK0rZTKcaUPJaDp5By4MHgqXykDEeT3lAKMnyPjlsaB3jDWrdg9V7ndQuwxZg
momItK33dftzwOj2jvgiy+17H7+33QBfz8dz/+cJlRshTUyLq+WIkRxE22YKKg/fwjztX7qW8rEw
GZwu5rcP5ehDlO0uukz/+v00W7zLxX2XoGABD3+FffQIt4wnFbsmfV9ZjObqUwIc6+NCzMpKwcxz
EaEgcNiJsmm0ND3xndxkwBY0Fe7iJ+9pDfVQhNGVWsabzSjuHulpwJyhEl6+7pA7EzYc5eodw5Oa
mygaFtxavc/DynvfZrK8Gf6b0+Lugd1uhTTcZdHv1X2ALyN4Wh0SeYmO8OY+lk4u6Wv0UOQbekxF
pfLv/ozImxh7re9Ltf5C30KXaCEkmln0/F7EbWJ+BMUKuWDr5OddpzjbKQwBpfWdur0sgUeMuRhX
6KdMfN9Tit3uKVq6IKCg8iDj+I4ifF2/m4KOPbFMwcCTylXEdm1TCaBSyU1VJLiEF6MjF1Fi6KyU
ohPIWTppVs2n2Gk6VhckkiPceRZo41mA4H425Yx3RgNca4BbXAHkSa96L3wEpX9NcxIywD6ZeM1T
6Y5wE5PFrjwlTkJrHiu2odv+exBHeLW4X0M5nNGxO3T+QERDoypzMXvmwJAYtMf9hoxbP/LE8+Ms
VzuP3viDdBKECWTtzTGSlJEfP+YNM3JWVif/dry+EaMX4j3ANpLngcwdaN50t27PTVBZCy/qWDCd
x2RTzW9mNV+Kpz37U5g8US0e0X0vaWpHmWg+2WG+3SuleNeHSLtBMEXK2XyWIK9FpMgXusHVdXsA
2135uQ+ATM8yLdNrQ0gthoahD1dksm9NLXMj6b9fWvUOOWUgrJCkHULQnwNIYARV9sD7mYYAiAsp
UB41PKSoRfqUbRVHY/evxN5soTHa4hFfSQ2aR1YsZe9+YMMmBM3NJVGl8/08p3GHe96DQ6bBYZex
mRJ4xj5H3wAFh/yYU2Hk9rj7RnDdbyUuLmxpW9wfqnq2ZFPNWJNYdg1LHPdfIYzTRVT0XPGo7t5H
xiur17sfJtxPYRg9tyPuVrCEy06QfqCZ9WqdKzfh7OxMHZqqciWkVGX9BrcpZnSj98uft8cLJ+kD
bb0NBXxtk2NLPUeFKXmNz3wJtolWvMZ1GC/x8qE5CnbhxEGhI49Y0t7da0+Jg5XRT75EQqoRMqpg
yr9YcM/cuIgbRGiZCCFh/Z7xX8UFfirNRM5ZpZxiQDPzg+S7MjJADMoWIE7u9VyuaU7BvrlDj3gz
KHPRif7tCrB6ETTuSZWoLpN8NAJEbLurgM7CJjOb4LRRPNqi2bg1VEEn8THigK+zKPzwBMetpQkS
dMYF2fUNWHnVLTuwDF3VXaD1SFWFs5cWiFoadtmqm2LoaQqjueurVUVTTvnLLl0zAITI+UiMdYi5
NzZ/37uzRx20o6/693Mgr2BRUsw0pFM9avdSixpGunC2U5MNRPiKZq9P/gDUGxHoraLZUK/BWlet
9pCYx//9O+ldQPzxmXW2kp+XTkMN3v9l3NADAcaX3mQzyC8sLr4GvBpc+6d+kF9fDcn78/YMbOaG
6eGEmKy6bFfxMi7dOqhI3AukqvUG13FoFj6QuKjJgIZHaM+LsAfHL8InWQlWhIExBxf5T9TPKPP0
2KHX5ftkez4X8IsksddC4BYAYFZ2aC1qXG4I1bl30oeeDwzJ2wge4Tewsta+OOtpoZt8OsRKasJP
BoK1J+ctNe054WZ0+83XCELf99/ZjupKpSpSi/5Bi7icvLViqAd2nxPsRiS/MLdjtlBcZvZNxY7c
bcw1ughtWtwK1GilgzC85mJoh95Y3a6Z+tY/5BSPM9HOgQTgcdRV1OeVk6bgO3fBFY42IzCbh9bO
NuDRMgrBNK+xIztt+MDXrv/SjRauNyUlyJzjW+bQ9a5amjo5ZHkvIGkwGUpW36bYqlP4+y36GjTc
/A0OyD2gQ4pLrh0n97HJknUp6jNeN3WsZVyuuT7zatBEigC27FacQ0HFOarNehmbZuLrzvzI1yWC
tnoX8gx0xV7zk+NalxTz7COsFomuqy0BDPwTTgiQUooZmJtw0q/ErpZoJ82fZnNVChJG0ti5H+4N
eAhLmNg1t/mWebjAW6J066xnqY9y3qVx2xwsOk+yYh3maTtJ+wxnQydaAtw+qSG88dajUkUqY53I
z7Il9RPOpd1hE/YI2oUjnAoqqlUepTzpkFdP0IMVrE1Z/wPJFw59d/VXkaVHV2uz8l2g/NgnQVkC
HiPPncllDzQrGoQKZlNZaflI/H/lhevNf+urCDZcLonHOnVwRIcMI8IFGW/m9UgxWNVyUaPLtidU
vHOVM96maOaDOloXgMmQSn+1qnieQ1nLtq1+bLG/lACYZgEnMwrUnZbhK0wHEb4jX44I7C7OZxh0
OKn9++QQCnHtm7CZ0MIA0pUfJTO8UWUYL6Qg8YpwDIUM9Z+fW5gTg/YMehndzd5Ha1TBdWqUZBsy
YMZI6M5hjdteyJ29MiIzT7AJn3HYE3uAuyW8+ePJDP7GIfMkWMQdCcgOW12LWbYYyzKlx6RLjc+c
RX+CBEg14AN9ZGlYQYP6fs8awcvLS7PUmvI6/nW8m15lCZfPJZBEaDbOhu2q3zZctWeNTYFS/e3k
zbEpQDR11BPALADsNjFPLvwaSMObnGPBAUjIhIry+yn1ZzjWBDBjN2NRONZDW8XSH82w21Su/mh4
fPlPAIDjTMee8M9VPWlgdYbVqqQ5hyKQ+3s6NcgjZWbD6+TFVi4QRvJvmJabdR90wBTW/RvhMzOS
wwGGxc1n7Ep+YmJ1R6JYsPGDDYn8zyW6mpCPePNKMNwBRVnNAvskIiwDRTjpOlsoY3DrBMup4Q/w
22nTWRhMKwTEedtJuQVdUuyF2k0HwVONexnVv8dwvWWbKsJjX7njwuw9nwA7u6h7e07B+C4dTKDe
VgnuhFT7AzjiTB785J+wJzdUvyCYf5K8OOUsotJPVlouVKFBRQWFnJE2l1segK895LjKwcr+c6bp
PQPlQa+iYyywE4MxuN2TH7znzA1BlraSEqwrubFxFh++xKLd9Sj+TmxOQTBhBrornKM8sTMFnAwU
XsvVY875w5ubandmzkYm5MAfbqxfRR0zqSRyQQSAM19ucTP5DwBTU3sh+BXxOxPghjVI83kQeSCg
GQg9mgD/UWF4lDsK3+ahqkdqz3hXtCfayudK4+9QsQYEDKgpSRdf/Ezqj+JKvthyXqeCIQDaW6G5
pnZr/hrwtO8fWcN/dYUp2YCi4HpL5DTaL2b4wbCX7VlgMgAgSTYIQbNGClEinH9g7PXt4gb2+RC+
wk/zKWxQ5t40d/E8Ow5XGUCCmwQgz9Q+iGiSxpP8oy4r1Ca5FNKRdvh7pRl7HfRlugTG1xH2cBIn
eks1ePEc0+SrUG4IXP5/IhaevgVd4TE2VCQ50zgtryKuB65r1xyWKQu0SpHL443IB4y0iV0ROJ7P
lIe5djD1iusgTzdOY8PNf0QeAbU3zzT06gFc+vP+2A2Ss02AP6VtQk7ff6KSoUKpGS4DxtE/WWqZ
j9ef5Rv1rPhTnhfIdy8oenfwj7mr2V+qRCnT2w+WyrdHl6mbcqj4qUP1TuX+sHpxLW2OQP+mvqcN
fmk2TFW/J2tGoeP56XrIkLt6ir7tFekY8mmEmJARX4ry8DezTtQsBdXWoAVMLeUl2sNNVOM11aqp
5wuUVH8fJAra/eMjmnYfpC6uQ/fpDp0lBut7VtFXhnzPrq32jBTm5TEQxJePNmt0+ILFgO+uxRYJ
PU7L1Xy+6fzIGR4+etTZjKesyjPNHuGtlgLfXDxRCo/HLqaqwbjbANHWK8+c9JXMWO58g76jarKc
DKakkk5BUgh8wqIFjKLwlDtgR/QGbecg5oiObLgJVwEUDvzGLbAZAkARcrznZblxqAEbcw0KcGP0
eZv8jUygzd7hk7FTjB7iNH/yz1t+/9gPg0ElaMvMPO15lIp2mXJznCoQiGF/634w7lZbgqsJkkbt
PSYCKfuCe/Dp1TfO8fR6xztFafXeRRXdJa/8iM9bzuyL8Z6UCeK+a+CnVrd15hbLuM9zPFyQ/auI
MF3le+DqG0fhtaiResVqv0dXzP8IKld1o3LfXNLNpLn8yX/I6rin7x5RgPHgWT9+d/yfWly7Hlio
zF0trsjeBEZbbkHlKSufIoFgm2sRVFjdSC8BfsgxkxeHBVqjSdctZTrC7vZqleRUkA20o+OrOwT5
1Uxj50BprjwBLlY8YH1R/8w6vapHGMh7/StAFP5+j/6VUzlTaIXccii+Rg95ogyjOmwaubfgheQF
p29Ri8GB0Ltjb8BWOHxXP3HBza7WVItoecTlQvfBF8mgSKjXtDCptUxz5K/AaCtNxitQtHJ8B9H/
dX1mu3R/3cQpwWT7K+iqw5hPkSzdgtaWuPY1J6RFGrxVSyaP+aIWxUmqKNV8bT1vh4k8NV0pnVLm
gvDoaEubK/A2jJTUnv8s0MhhjcVqiIURbJhlH6mQhKcHn6AraMTj/8eChVOOH8ht20FRSUVBY7r+
Yujy2FjHdh6xNOq91MjlVgC9ajSIhACHNiJPeyX8FASMmfHlA50UnhxqzMMB/DSE8p+auUk8mur0
ZF6KEuAlIGAlBuX81TS44rAt+NGVNDoVtANOJiZQZ1JNCnOfUB83wQRbom9jHFaxkIpogM5vl7+Q
TvAThpPniX8jiUerrUowqlJA2U9T3RtKAR/NHeWPS3u9om+832Q4flHDjEIHIUO0fQZNZMLSp31i
XcwRCCbdR6P3o8H7KyAHy8+yMBoIk49OoD5D3/OYXbO5ND4g8xemvHi3LR9FHxxIUEmrGCmWb7na
gFmHipz21Ie+PSGwvzYN7WCyhyFIRTVQhE9zsqlVuKIKAP4A0lhTO0skyYGZFGJDoaEKWKJbWIyZ
k7myLhpKH5oBlmZ9EBfHsmAMDHaFbZ5TnarEBVt7OKchoGNSCtrrZakkhrNIT4sZ6MNWeLmafREr
YNW3+iQcgioLZn+ketu/F0qOmfrWcXdYvShoVswzuRES52IASyhkQIa5W8sxq4c/vXeIAb6lO1N7
D6gjR3JawRHCLPEWSquNbqnfbJYoHSIDiBAtFGJloNGOoYmfR37037iObo4zdc/c2CVcR/HeTv97
oRiNIr4dSW5X6VEOUd9CN4wPTcxwThGY1W7AUggeEqEktJOe9woxYWnpjcVN8ONVNQzqr0H/tZ+Q
SpRwqkUkGP2AX99dFJvEEe0CYiR7FVkzyxmjC5L+LKF4lPWEazTiv1/1OI2dGhYBuHLDvXc61mvp
947QG2zNrBywEKQ1ReMWdkr8Vqoae5uvyBzN51Wd8INfFAyUErWSFGuKXDdd8YskRMaK6gEDOb+9
2oG7bRzex2m/2GKnvVxKyVugr0OwtxjRtDW7KrZ7eGKMay1HE+uKbwlyI5BPTJM8qule6wIohvg0
suP+V/XzNWO46kz9jy5A8ZdJIkP76Xk77OhYBVWZIfVELtIW/aH1xeXeWzpnm5yXlgadmip2tBld
E23QzNy7JJgKesS7M6g/k3pITWuy8Uwxym9W4sPMqtdvtRM0ZbQke5KBK7zKRqXKo1ayRcePblRz
4KlTOpPCCKtMds/QDm0ZKoiOUWDC8cjymFVR708ZkkFy/Ma3aU9i8aufg4TN5qbv/h6aiW1uLv4s
/89M5/nJgHUy3iMaacjQSIDK8ykrBFsjyjeqAOrZfpuPTTSeV3ECBpppA2XxMGB+hAzBVd+xydmC
LTk2NokmFeH5W0Ccdae5kWSYgb9H//y/kBlYu9J3jx9Ls9hd0yPNbQU79sLB85tGsKCT7lhzXDth
liTe0bv8NgcRa92obkfEmdRsnvTDbgdtEnUP6TxOojvZBHSr9URXDhyv0Y9Cd+P0L8iflNAU4s4J
qi/LPxB7uinu9TCOMURKKAXOQpe6e9vwEhZIrbbvcWAnzNvcfl66AOrOtp3GZyzVsaXvhL6+Xbvt
lrQiNpMbMADPWNOgpAdMYjvAMPHJMIz8KOyliZI4gxVcVXiLUVRBkj8/kGzOX3j/9XiuaMmaAqsC
qpIwuw0vNgOXTOsi7r+0COvXkj8plGpmZwLlNDiGQk/QmUE7UsAoYM7sHke20V6Qv0XJPpBZrXzt
ntKgPTX+F4RPnB4rp9BujSYRtCcVybk60sg8HaQdRJK5dUHwPNl6yQqSevxvFn4bg6dfON/whRRV
//qIJ0gapXvfPRkHbkHDpW952EDVIk6diCTgxfyZ8ClYv9ZtvHaEu09WBRs6CZAnTrV2qIFu24r1
u97+SrOeqyFSDWd/adcvNe7Ri7d4sRTBhx40OlWcxtuXhqqnw6zUK8UB+YXqQ1WbcmhOxmQIkI7m
BpIi9hmSpvuz+n2trm63V+uvefV6uDaPc9TnjkKXJWPvnSmjte/F30q/+giQIk4CBjGFqqK9mpLm
Ssoj8H+WLmkYK7gRW72sqOcI5z7dCEnZjxjTk6Ml0iMC248VzW5TUSmMcO8pMQeRHfDsxVnPfg0Z
NbJMzbfmZVH7Lx++4mkpH4n0GbMU2tydZEwW3zyoNj3gzvsvSOeh1yndRiyVBbAnASQSrrkYoYLS
CgQ3NUEENeJrTyQYEr6jTWgdvYluH5VJJc16W6qBUzJ8q0mO0ZFfDk6Dky371I9S7lmMcKtUvZa5
nTNh7GlmuT2e5jvcGXUYd+B05S657YXcSZCQWe7Lv/HzcvHVN2SXPNLxWK/LpWE1f9KYvjZpK1kR
wV8J0IpXNQquINSI3BRO6MLyf5ENEXWOpXac6yEXj+ZklQ5GlJmlN/HyKV4DOmUS44gO9wZ1ocP5
AJF2gwuGS6o0dFDIT6QD4CdQo5ONgBENptqF2gAFsmSXOlvth3kyGYZPTiWiX+HR++taU3n2NIh6
3uokWJFZoQfrXVtPLPUmOebQZiA2AF33IL94zQ1GKoFnZbhpyg9S8ibX1bDevAIgxVejIb6Q4q/u
DfhltbRAg4gC6hY91g5tEGEImj2mRCRTx29un41JlD/jnOOpUtTn0HXduADeTTViT4M0QsRgcsb4
w0n3xa5gA0qZykZtnG/ZZZa/pVbL8LAbWXtNfCkwBbkLcvOXFxBFlGq+q7BJwLVi6OjnoPsh8VWJ
Sj49fUSvcJRB3EoFekjeaDaJEJeYAtE+rUCPONyYk2jaI+dBfIeEMkTN+1ATVjRxPPEC/hA0yWnj
TNVdujzmA0hhhBoLcP3WzmOOWIUx1QOmir5x3X0Bat53TEYF3oQ8zJ5but2a3ThmnYkxNMvQZ/hF
VdXPk2dXPHKuf1Mc4wIrV0YBLbSmCOuLub8qr5TAcGF6yyYeiPtWyM+wfwGnBnBl90ti+M471v7d
pDlyIO7clexBN6e7tdDeuSKTuXUvcPfU0OUgWyaB84XFzaSD+5lrKwbs28Opk/hXozObOTPcMKiX
mJQBZfSb3KrbT2us6WZHSc3OzOyNCVqGqYRHqJoNnDgdVi4dPWKrCFx+c3MLRJKn+vKGrmsHIIZj
bpZsln0FXIzfV0xT9X2p5Ul/ZijAvHl5e8aSQGF3g79xpxBUjyYG7kBBrp86AGFzQVi5f7zKETt0
sbmkjp/qFIktUeHi+ez88wIUhDh7xa4yEzZcD59j9dYOs7Z4KVm055NZPBhzDPDow48PBjVDffLX
UmrEvPdYXZOT4fvOVBU0v3dYrhbFm5nIJ4r6+dfz01AARKkbBTan4ejuslBUSIsYVoFZxUYIPlcq
yJW5I/9kbpQ91xjjChbgz59qnZ2jucY/R4jXXg74Xx/thuvQFGckEjMfpENTuhI+t2MsJD7E+wwb
fwKat9Jry9SmuesnolXDKanSQmECeFJRGT7QAXd397hgUAp3zn0qRhH+PEFIDqJ1471fMy+Xkt/t
vLF3w2nk5tDKcWb9S0pUyLCyJQu4L2tuBmuCrQiF4t5dHYxyCPTb2+ftdncJJJmHtKCelrbNuqvV
pzCEJJ+yC6TQy//E2n4ThMMgaZMJetVnN/F+HhD1602oigKMA7A2p9Dl8cxiT9uZg/qK+9KRWuuG
6q0NfMy7A4KIBXU04ug+m6hbpM4wosKokf4f0OKVV2GbYYI6Ikv91UZqCnSLFPJXm5JtWqEBCOiU
QPZLxtbK0fHStIRFONEJhldRl4K5LqMfUAVbHdP4zhqtmyU6VlnY1yCsc3TgODAUvTOKrSHKesVO
99OJu7jJYstTTerxNXt+EAjbAwijMUTUMTwXYZLZep6O4ENFrGLyUVjdQ1t1E313XNVpZHKw+0DT
yT6oRMmaXUYND51qu9+oLfgiix3oq4QENd6jXeJd+BNM0Pmvzob+kJYhNmQ/NRxUC23fW9C+Z+VP
xXlPIeDy2Im9J0vTqzarGbyheSUWzLLGQThNTxL942plpsxQX93nQkmXwClRqsrFNaevyiKRw3Q7
4qM9YR3TIby/RjN2wppio9o2HTI8yECYKuFmHq9G07Stcj8CMhZotnxguqHrp+PBAUyusszTas+u
89k/8Y4IgVHU9KEhxpl8F1VDDebmvf+v49++RTrgC70dWL/j4eZH6xoP083NFfgipAtRY1iQs4Lk
gA9x2FX/NcXQ/wd5jFe7Xr5NuWhgmZmalWH2Y+Y9V73xxGiULf2BvDwt6Ziq1tD7Tto11pmJJ+N3
3hnMReXQdiXVvaQdHQ5N+LeO5wApybk7HMyY+frrORUYH+HE+hTpAAiufMmjVGMt2+FNju04kvif
LL9BZ+jfHAbpAmRJT3Jqyw7JyG4s2n2tmXW6rxg+S0Td88V0LbG4UiN+zEh3xu8K3J46Q/4W3wJO
jlGuM71TUHXaNO2nLkdk2w/KDV3mWBeqZDpkTzLwPMlyXxAaJvZxWTI4s9dnbgZh3qYti3ASwkH6
J5NZ8MG2ZErWa4/bgF5cW3GfII15F67S83oC1+ydRM0djokjDOEJ070ycyf0G3GjgYGDUsWQz1yw
9wb/uiFpu9uFD7OGe4EMSn3B4+vuGvveJK12gPZVMHAP2377VRp4/DSF2ZRV/msHEbTIgH+cG0el
PruxeQRf9mUIev/vrN4Z8ya0MgWn/FD8sJj+TYi5z08P2IsV6sV4KTIQWKOKkYosPxrn+7AT3hVv
2aFO0fqLyeJ2PI3NgO5ct79G3gWGR4BRfm3Mlu7SX7QaDFze7metlD/EQZII0M4J9h+JcmX/VvuH
7ua5xfTOLNufUld2FBM/EcYAYyC8+kXajgVIgWNtXZ6okXtOGl0Ub9by8ZRacjKEHHPzuYjYbOlH
jBvAsDELt5v2/x84U+3Rni8Xnrt1Q3nhHeDTIW4KQKHOzuox9gd9CDYeYfy5eeMSBAmKYMtWEsb7
x21yOxXX7J8w0vHQdDp/5f+80nlPeyjCdExfUP1TvE90S+kUYleWZUWWe3vmjrQCJ+mhSfB63ish
7mcXVLbXDvKysQyv5JraguuNAUSk79Cq2llYiCE2NmeAeKRdk4ICyXZN6aL+EplC1pEjgtbHI7Sg
VnW6nw10JUqM5xyFYOVrKgJ+taxXIjcAfml6EgqfAHZTJOfKvzQNuB6yczjHKtyUiAgTyulAWAeM
Z8vyTeZt03NbclhSfVeshC+vHj0hGbRLU5fYg3doa9m06C87pBGLhPv32lpyh7ZOk3IHDd7Tag86
1mPffg==
`protect end_protected
