`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
fjFb11PCHySA0iDCmbnt0Uu5TahbB0n4HAlQM4dSqm5Jj1f1u3O4zhgR6PNMkjWCudNh5jc+V248
J/1nH211NA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Mg4oysUv/jIIaSb8YNti1CGwNP4sfPEF6O726w2scoYS9ZfhV+XJzhJFor6p1bfQR0J84gq9SSJe
cBcSvsg+k9b0HqXnh7netTM5Ure28p7uQleRz757VYh2J/EzUDeV9eaP8Aj2SZy2pRw/6FnlIUUU
Up7tEnerkhln4SdT+Mo=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
Ji2XWzr9x5xfAv7+3i8XDINnXxzAxFJ3OTYREmIQRVwJFyoPQj7JOVZoOAchhI/2ZCyh7oMZHYPr
8Bdsh3ftu1jyAOF/rjPQ4vEMLueZ/FJqMzQOcnA/6lugsrmlCMV2jJivfnRV426+6oDXradGMqOZ
1dlVjDlIiqhzKaQq/nw=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
zS7H20N1boSFCvzwPRMa4J859ieSVjyRLpF1Xyd1px3elAg0zvTYsPUWxQ5nAablDb/QhtKkQMNv
0fuVCn8QHOeiVWjQ099l6V96Hc3KjmiZmbLX81S3QF5WPlbcwGRLDNr8cgXbPRnwRCcMW0b4IxUQ
D/XfWhnvHRB8Afmi6TrlqhBQcxxDkXwTwq+snwwJ2tTqx4TvYUpwvxxdyknNNoYCZR0CgZerBdX6
KewuxV33CqnFbB7XUzdJFv0FkM4imN1z7KW/614al1q73LSswhk5TGHqj1UUdlv5OgRGwPY3Ke4L
ndz8LaoE5dVHZSZpye1mncIzYDV6W4LaWGStwQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gz8KjTYHavfCWIfxV/5do3RS0W6z0r1S55GzScyTAEERTMOa18giEob/2HqkDNWrWIItAYxnUWXO
D7qVS7lRsC0C28Hpgw9aZ9+73tMtTzrGfQgCZhTTGbFv9pu8m8HHa0P+TwSPix7T+sIpGE1UVxk+
hjmsUPgw+qgRYviqjczmqnNP58iVm/sag0nO88Izkr3UFmWww3Qu/xZUf0dl1r+jyaZ6OZOfKfYk
HiCquIjnth89hSZOHE/FbVaUJ+r+gAMC0SI2FrFZEhy0+eKqZQBW0baOl53Whft+a8sgKh/s2rPh
ZH1RF+fMkVeWB5nEalotTGxIGkmzuHugRXAWVg==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
bxrNF2OuH8aKUy+g7Op3+NDJlme1h2O1mmA1GsrEV2CnIGOLnSZQNDPp+zT3N7rn0kbUlmqcY0Dk
DwrLJ8k02oaX0F1/e6UgYluwNwByuhip2tuLRMaosh7DjUrfHenA4/69szDs105Mit3ZIRt7KUTd
JnOEUnQV1QCLUarV2Ov20s2tT6FBH6kz+x5s/39edp3HYJHOVwBQ5PM0gAUOKDxEVJ07sT46zDGC
8KYJBQ2mt1dWvsGNP5STuynUnSLahhLaCN0v/7KkH0U6FzZUGOhQ9nA9/chrSJG8jjtUgHkZhCXD
zagkLih2Fjb8mZu4NPweboqqS2VyyTbEKHKGvQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 55424)
`protect data_block
MCURu+qpPjwTMV3apKdjx6vwphvlNcjoxjZV2ZjfUEP9Qo3Gb0kSWRN5O91MbrqoLPj1X8TVWpMv
IWnP71EVbtqsE1S2ntzIKXnO/POvA6lFY5R0KBQ5mqwUHaTA3BjxfFpj219v8fFN1VWGmTDwb2EU
9F3FFxaVEL3c3ilxl8awWxZR2TUNp/QTNskKv7NRdBuuc17Lu4mdMuD11k4Y2ZKlVkAkEiPvmFbG
Y8ZP1P6pkijJXT9byGDB3/Lqv5wqyJtW2rReJmeycg4af0K1BmBVUtJFPMvrBEKBBkMK/PWBA5Mt
E/mSuwgCZcO8wAfKc77Ej7ppFHum5bpTm1AFHAB8MS2LQ8zmEWHx7oKbnghGbnBMk6DFkavcKDCY
Mp+DOGm9LWEb1S2OF6pAN8w9O0gyESomrmbtclJfKJawWRS91bX7MNNDaKOpNR6krhLdO6X8w4lf
i+aCPHLIcpBjdAV9WMFkv3HRcAzkEUsOo+yyl7hlbvF9NORZ55yk9FdLEdXn9c92PLD84gRsxrYh
u5otqd5UdE3xtjSaGFfRtmV6IG2/K2Kh6tHYx4e7Xu2KoK71J/EiMUBGf5xU3AlTSc5txxoF+ZrF
PilucOtaMfD8qk3e+8JYs7dykGSefruOng+zZ1oWZWtlieaZ14hhkI0quTVURUGGLHtvt+BhOhdW
ndMDCirqtSYH/xDAyK7j8VhmymPF9U6Psv+7AHSDYdBRYkx+40KmjO7Zn60UQfozY8JNQE/UtfBE
N+i8udXSOKAUWWlAtzroTlltLaHqFifrKnuld8b0T6uVS3tLv+Wj8LkhlO21GjWJWAj7bd9kSBXH
ddtbeqq00/yW+GI915ml3lL4YwFOQjMDucaE3xZ9YV4OEZDk69s9RSgvC9A5Nf2PdQXr+LUbwNEj
lLPiwy/vGIEfli3KY42jfMYTgjhmZknpoAU8td4lUvD59iRryjliZTAlYSKUkVmuMdQ8BnfWOS14
5TxAMOO8Ox4a85m43Jw3Sq3zUvGYqQAjxWqaYheqeEER96/y/+ZsbcUZ9Fw66sdDR+WuLeqL28V2
q+CtR8ca03OPphMv28gYL8AMcfIJ5La+VDxg+v/2cXN4XYGVyx12smE45dYxC3/NsI3LajBsC4rH
di/wNnM3T2Z4CdCeG1oP/K+/KThVWuGTGMUvISV+JSDe2V2h3diPUJ4JTS36BF1akPumzPino5RS
cVG+iYBsCOXR1sF2IRm/Y8+0s/E8Q0X2ONE60bxPdFEsXU9s3oyofuKGRpDzbAQXQ9CigeaFrDgC
zVlUNPG7t9q0W0vEPxlW+kEkTKW4vq2YaF+MEguyWbMh7NZlIe2QtQnYctK7CCDNHLoru63nPEYg
14hFXQZl4KsmN/zk2VVWMOPADRSuzVfqfWbcnmdsGPjR0tjKHGyjCGTJl5H53BRYgvum6vzXtIa0
E3Zq2gZYOyOxUF8Yt+pMfJm3qzWRPXtXW0Rp11hcOff9okiXSpZNogtZAqaBhHV1bh7srwk4F/Jz
q1Dxr4GsASAOnF4zJwpKYasImkVPkFaE7UxEDHld1S3Zb+wTJEf0RlmMpt2Y/ouH5upxXnLfD17Y
peSbaE16wi6mxU1tFrTIVQTxLdEu57qv4eWkjqNtv3RjL+ObzYfDyDRCBlK3jocnw4dr7lSV/kvW
Hx8v8MuRU8F2nV9glD/Efhd+Ky5yu6Q7rDA/U2JHSz1687G7M8YdMtt7KDIAqQawzuIfqBu0a7r1
FZLKubVO07Jq6rxXK2l4HK7JEHYqPBQTe+HERt+qLcmFzZbWMT8HsxF06yD5O50FMyj9DEE3CgwP
4TBAVVjFOHYwFsdpy+L/67habf3Kmj2yoyo+0M/BwXfOEQ/WCgyh0fZ7m1o+pir5XyNOhRmpucJR
NSgumVGcyYNxU6XpYrYDNK/jQCfvvZafn8BIrO/NRiXFUCkGoGF0UPbDqAc+VbysHXHPGSGicCee
8/K9LTeLa/p8IEoiLnD8pLqwJEKi9Me1zNsI0oit666r8s7S2IfAwJYkIqQXH/WiQgSTPZdMTy+u
lbNcIyF19vxSPBnIbG7IXv7qaXFBFVfNO+S+Qx7ZkYJMRw9adwfluiopZAeZZCku0jwmaXhg904j
ONcI+4Lb+U463HfSa1yvQHZnRKlQLgv0FHaX+6wTNADiOLGmkpjBo/Lfs3mV4rvb+DtokluEF/IQ
1WczAX9ztVCty0uEh5V3B5H1rnQ9aalkpp8AYnOBkQmaArOhtakyL4cVbYm9IC+VCan1sHdl9ZhV
cpv1KGcWlw2lVsWxldDVGM5AEuCj8sjfBSAbHoiUlBkeNzXDtkc0jSEOcusekEHwzgdrcUv5PzpS
GXPuFvaliIscW1/lqFaIrMVOHFF1XUGAh8IbnRPYuhwTNsBYDGwBVRtoUI/vVFI7/YFxY1QxT+0M
8eA4gRTsnx2LKLXdR1i59rT0zPjUupH673rZPnOGdBfsBIrSvEzCOGbo3yX15ARvSTc5Oo3X/Fpd
I39RYM8bWoDDPzDWNoO/8u4VNwvPOPp3tEc+JUxYt8Brf6rEzSDHcid2AswL+uPdUA9sMaSYeWbz
a/IRRGCJM7o0BAtDapQ42IoJ8B5hta9gsIdwHGNMzcaLxnhyGMWEfX9adySNDS2wzyjkb+n1p1GN
DztX5xAX/ZIYvrz46JJTpOxtW5lFGDnwL2mwmMlte1lKHjZ9eNNzBPd1QhCa8LvEYTuqR9wLi5We
2XwitGs3O8bzzbNHQLnh8atwcTNvwiM+yE7VwCiuKgGEId2jf7C1yXJcEoGdbs4gu/+565gO5rnw
USh+lrrZoBZ9pe6gImSulDEVKyHgT13EZoV3qfLZfG5HnWNV/mMcwPUuOIgxgxYqlxsBZ33gaa2F
k9LOovu42X+vdY0gpin5aicDQ7H2Hz7M5sac+/F8gwa2bziZxmvc2/cUdWP5xPBPin4L9fpEAgf6
r6ZQ9oMzsJQO/nfJwvhLu/PmvftWb96hrLwqxJ5qhIb2Nfub3GntHZJjRksp+Ca9OtJpsUzteW2C
LsPcLqjUh2R7kZyloFXK9YrVZIN5P/8acbau1+3Izu5jM8x5uMY2h0QD1Kd8XXxPH8UvIhRQWTyg
vHR2mj8M1H761LnQbOyP8gfH9TqXGwqXS8TVOUxuTaog5xXqKmwcosACWYXLpEkUHd+LJEsFdD4B
Ewb7S5S0KcnAwa3bgEJ0P64s1gOarVa83WxYhWGfQ0t7zBHf8dId03CsGipn2zChJ4QK4bt96vTN
s/Pjtx8oRovyFc/qXZjudYgr6J0q+o5VV2id5RldKJq//HOjusBeigVNTCfvDysxdbwW0s0SZtLJ
4lM6Fg06p0H3rG0tKVn4sk0+6skoGFOuXgriUjnKeLUSQPqxsmD8hrjKZpm1MeOi1ueRjUJ7w+Y1
1obSXoppVa5pniLVrYguhn47V9E3aN4GYX+2cpBE6hcPtt7wgwtBp2xK8iB7JzX5cqzXqNkhCLSB
3EIkLMBnqzNoznlZLv/QtdOoXQ7d1gY2VmW6sbsiaeT5CnIbTKWK32l9Z9w/ZgRtfdlV6CkLOWYI
g+G0NVTGDgzPHHg6XCZ3dLYOKrZ5dImvSPXxvnpNuc4bnTV1c1Ueg6u3AKvYXdnjc7V9M7eNYxb7
6B9Y1qy14fQJPYn8rGVCcaWbWNzcUmt4oJmvO8YyzD93wfSIt//Z9FSO2FfVoTPubFaMLkoO2kI0
ny/smC6filP3pKwD4GVaCONCOXz8a8pOGmgVOr26WNih4HvjWQxV0QlVt6VMEooyXB3Fh/AVt0KT
gR3nAaul5F8W6sCoNaX58BdD9GzUZKxrlQcyngBg5k7jOR+NZ2eMs4klyvSWAe8rTbQbi9k9WRHo
QSjlzcEDYhtTLhXwIuo8AT7T+cSL+P7lV08U+YleFlfptK5XHWUvohtUDVeS2+NPtZmAc+0l6YkT
ngIgitjXIjg1mdT1WlCpU0yezqQfylVn6EBZn6xoJVJGgP0mb5cYWGOjD7+4iLNMRFnCaydKM9K1
m6eI1uyQ8UyeNqDEyF/nal/G+xx1aoSY2fXX22xLex/lkuqlznrMJ4s2KsSho80/XG/i3fy8cZyH
fXAuAc8BAaapZnRr/oCWNmKU6gb3Huph3IgO8XFLdpWhAmtuduPMdSDV80lgbyC57+zo92L9FYDb
EcQ1nDqu+2W3OAW424/yxtvKSr4QOjLocrbah2z4mJXKpjrIfJ89QPWlJPUC8Nj1ynn7IW5vanG3
VMkb2FYhSlbXqN9CRDCNyRdM5o5hTszbdnudQN1mFsApDXnlBSNJV54ctb1+2X+5J1cgfAxf1Guk
mLAiAmVTbYdtA08OExbca7M6ytsyfLniFL3isuayWvtJDd0eohzxHtF2/9xWkxkefBOcHdttXHny
VYNqNZ/SykklUIQL0uHWd4KTzxnZTED3HmhyujoQAxgRU9Pb50Q32JjaEEmQZbfCVyVFbutfKHLR
4fpcv1/R8ftdtUfUjnJN31v/JMYeZlaHOLmddfwoedU1JKMATJ/8D/bqq09K0fnOaI85KYmmd9u+
9JGYIUetu+zR3KAswO4u8ax+kIxg0mn9P+/n9bFkBrndx+6taMLIZUGxzq6thmeWgeRhSdOZRW1V
WJC7CsU9mx0T+AiG4Alr6ZLrXi3mPp5g3MRBnn01YjkfzNtBH+gVhG5q4NL5Sgxbt6aa30HfhhRL
TcOlstpgjhPebGlhHlcTHQJSv7EVOY5reP5FAMEI51mk1uBFN/Nk7r74KDsYc2tk7FptSNFCpRP4
f7iBhhlht52dSB26FeGeNZs5y0rtCIDdnVneJwsFjlAqtVTYV1R9jvYdGDP8nd/tDjvY9r0voEaL
Ims1StJdELETCDVT6uj7wSl/aE9lq4tMA+5iyPcw1IJqS6a6RWPQGchYqb0OHwiybm00a7jCzGk3
LEp9Do/FZjRrF6U9UaVLllAuAv3inIcXnr0QmoBzUj3gIN565KoAigVZ8DfLg2TGGpOFKJiLxtvC
rG9r9255OTqjI7obeQhsuhX55BbQdhSvXiVBmYzwkOFto/qp972EYx2DLxKzuqeteClLP6Q/AFJ6
1kDmf/xBOg03c7CDASj6uSipr+GEvGiy0rOUeAa4IiJvvb8C5yc0G2SwjVChN5//PiefavN0SQrp
IEEuAVmKyfxyWsq2ZdjhnehNMs8yuPhOoZYZ7jCQxGs+Fh/MEtrJXkl+k9sfvIO35izXCzbRY8Yb
2wYNTtVRYfgxzHkk6WK4ufIbi/uBkJLptSJmYN6xVI2u6LuNfj86dFcdSrxMt03bJryNSJZpqgDV
OpckDhwEPIRyhYwGYrFDpfteAmV045oJuCdjtDbVe+IEtyolXmt2UTpettaANg6oeh7bXaNgNrkY
DlOkz/xEpfpw/rcwaGayTtySvhV0tWZaYi19qVWgPviHBKxTX1v5f6vHtshTtS9WaYznYVybYwYF
JlaZ72VlahUxIdd8amV2O9w31w4COqu0iBNEINUQ2/HLTPhaTem5GEzSi1uB+e0c48qm83CY8t8v
vkKn82qjVJE9ZlBSWMZ22PYoZnaiIQLuM90eLh012YkB7cNad0d9eHcGAc2lfFN4/3PVkR9VShZj
Bf3vfhUEvx1t6rmMSaOl6k8pGzIHZshrOoN+ohVN8HHkpovj5aS/LcKCAhkhHLTztBgFOxuoZl1y
+W5Kaebz3afxS/gh7hQ62HvHpDokrka+AO10zJJam3Jsu6Qw+IAChbvjyPFawsLkI/G5qCqzJg5O
nu/EYZWR2x3LkZmFrG8M3nozNSJN2kc+GULMLUwsvkxj+CtvvZV6X7sT/ISeF4cLE5In6YA1zfjS
Xg5plNdxACx436mQD0tH6v+nupnXatQE967jILjgvyFClUjt80FGZDO4vieDWbeSF3wnn0yn+IgW
ainu7ZTp76uUaG/QhZZUumkc0ub5IDl7xyGjuy+OIxjT+XhCzlG/3oi3U2QUZvRuNvn5GCRXYUEx
07YLPwXWwezsmszDqh89zmSvSd7VmsTmwTusTPITR8GG1IWOo+tS7FZjSvR7x8HcvdEk6WKDVhUQ
BvVvhmDZIfi+lz0Ja0pwXI5Cc3LBrFYC/okXtMhnt7zTzEYiBBBo3KdWhh1RWw4x0dnylZtkIEE9
fqAefu4HVvu3O28Ig9Ss+4X/dhDk8er2Nce1PeKRhWpbLJ8/YIlYjP/8j+FLaBx0FLETdYJqNkdd
e+lWq0OtVCQqssFT/WInXHA35Zeivllzi/wiVM9GYg5X8Xh20LZTC9D19uH8GbKoo4hsnD0qd7/A
X6xsmrEf645unPMS8IsGxrXHxslpcpoCv+k6luNriCPGq5tdU9xNIA4ZD037gfThnRXt2fqmKeNH
Y3xTEwZnyzmo8O6SEvaRi3wIPX1LUs3fx+XCT6MnNJZoa1/kJUJNYui7QpNqJEAmLwT2xcuD4EKB
W0/fpvI8q60ccxfq+Iyrqpp4tj4JiUU1MZmwfPwqCSrkc2WyIZdZYVkbH+2uZ5ELiyBExr5zSokW
U2dcZb6XtZB4nSBGOsega9nGAGiiEgncZf3ML27i6r0MTWQyK9P+RGMPop2PY17Zm3KpuLQZEWA7
LAECc+UB2PBioLamH3YOA5udYeu2TZLx93nGSbzq6+A/TRX/Bk66LV4o3jSlrNqqsETlKhsWlKXb
/81IX6GNyDbD4JyE8k8sdurxQh90UoW3aA/v1s9Dc7X8bhxCMNYEvnhGAJySIiwAgrtmb0/8dlJX
RkrZ71aq/BP0U/a6f7W3fO6mknsW8y6WBVHJfKjhUagNxaz9rUKY3rakDz5Or7j4SSXcJrpB2Fft
1jgC6aW6dbp0szzVVCqptBQzxSlIOJedlbX64Azx8PnW4xWc1MyFb2ABZNyVXoqPu6pKWXbZrKEh
AigStyj2JItm+SQXa9r2dyPIE3DSPwRAajN/GeCEiaqzFRAT4L5r+G7cx7Z9Jb0tBfwKoYH00EVy
13wY4V/ATA5xxL1zMPGWNMjGK+VQQ79AJUpb4aVM/pnAafPrzh4936X+ggJdbhOr6aSyg15YzE2C
XR8mcwpOd9BEhBWW9NmJnwwuVCOqCbBh+7hzLbmSgKmFtDIS4m4GCSQQgNRfOxfJ9kUbqQQjyEgZ
WDvHtLuynrdbqqLegoxKoBHm2gqtzLJGuAfBUKDcrZE8oucLmyQn8HmHvIj3UzSKuhxs1LY4gRyT
NplmRD4teO3S59L+JK/pl4UFOccKwFKzKotxpPCY6yyMc8wdBrmSkap+uTElZDsDTA5jGAQHNpis
1vimlBIAif/9iaigoPp942ETYeRWHhuWHkAbRtssUAIgSoONATjkG9ugP2Mp4I5hiEPKJt2POe5S
P8J1xgYlTAJS3DqquLKP9Iv//kaG46QJhwpGCjNfKSNXLCOsuOnkr7tefLtFtZcL8U3Fr0ooLNb4
eIF3Ytr39+lBP7N3fHe3i2g6OQqys4uZQdTZ+B2jlNrM2SPfLvXPZuYEVhDTdH7gdq1yQ0tNDap7
5yVIrwgNb4LNke0adA8R82FsN3Qyhq83mBS12KDUwGBLbeWDgDQ26lu2xbZkCAsftdJVXkPYF1i7
SAvwHp8u+DoJwiueAAuofSzoj/ngpEgq0/jzMtuE3ghDIxXDAcvZR9MI+/P/tEXaOcvGxIwnIeVq
CR1SzrXPt3rM9VX8cuWefc+Xsvo+aqbHxQc6/UsCwH2ohPQcNmiPj4e/+m5+HngU9giDNAvhmsP2
lgoirk0kSRpSCbukLKT0uWXOg6vGANiLL9FEubV0kdkWfhNde+3NoKlZtURvhZEiNP4whW5HDZtT
Epb2rZu71bbRqQ4DkAvBCJveVurpu60Uss9ii42FCf10LOlT/a7ciucjb8/fH1UVPtSSccNzhfJL
Oqyk2PD+q6knALkCaKjaeRMJmvLKA25bWEM52mCxovpaY3Uhla/PL1SIrquworwwjVqPAfvI0uYN
mFAr+qZ5gq/4j06hMGY7K+kPT9N41UPwEHjtg7621tRn8jqYQ6gCUrwiUau4dpGVEV/JgtTR1p15
NrCkv+urD2qnwe/9ExsjsSBIYXAhMxbhnwb/i9uAMbxXoihmKHOOpI8IdBpC7/W6Oiy+YQe7AMH1
6VQ+FoeWPgTEg/gK2H7zLfCT8Gjh71FHDmSXAh1db/2bqGrDiUKNKW/UGohCvVAtnpZYBRGDv0db
ukQqrDhOTr2ZYCnj9Rf4p0Ru3/0XW0zvskx+KN5xiPR1Nu2XRdxiyOq6RmYw9fHWcKmoD4GLEWB6
CvS715W4GMDbzoS4e3luSrgaXLwtSuazhgjLfySE3L9juAb9WrYpIS9AWvIgYgM0GryJeIFm6qZU
sQWce/l3BQWkqtgEvSMXIwUsY8JacUmC+tNeWXwwft7oXZSJIwTakE1yfDboIzMzArbMUIM1TulU
McXDnNeab6S9YPvDvyjDzIydQgFRur06HJd9PHRXZxtXUZXi6ft2WZl/T25TvBz9YtDiQOHudJ4v
a/BeecFOfyLke3vPTc8kmnx/Udxp5G/LBbIIjg07sE1RLKnz7ImViawyQxX8MUtnyg0K9wxUklUK
WBR00teRSjbpG+UDlRfF21fMllH+bIax1nqLdmv8u1BPMMBd7BrXxLdp+2W/A73+DDOiIFpG+a/E
LUGtmXs8826K9/1YezoC0AOUBybKJdk3aAHKQBSegM1ahFyrMLDazmgvRHm8Hw5Aeqs05C232E0r
l0G0vYWQ2fHOb9xl/P0RzqxUq1s4G/YCmQ+/ePLJ1jx3pjCy71awesvXmkiZBYZCAqkNcHKDoUEo
FLh4B3GNCT2IQWcjE8YQHcJEz5QiMNNnSe5UckA93tH62yhUJHebYC23BfTG/DmeM8xqHo+QI3U/
MMC5bL5OW5SMr4njdGmTAYZsrnqYYlmp/4z7Ay3NcOJsxz/lZ1H+AUz4OlIyh6WDXI4wux6Xa0LS
/5mI/+szvgLHYzGQwN+gDlaFxYdYwLwqWiOOkeMZWEKqxUFhTeYyZxHPcynclJHEoi5wUqNFVxls
t2zlARhTy1HrZ/2UlCpDcXqhmQMwQXGWGZBn6jgR7XLDPoUQkH4RX5VljVSMNWyAY55RdDwnm1jv
nwlCT+o9kG0ltTsqjs7iBx74/Wp/rj9N4J/LaImOm9I+ir/0mTbzIhVWGbSGohPPXFXxSCa+uzc5
7sipTuONM4ySDtTjHARh/djNEUgqQRupKcgzuKIuH7wb9KwJ6lOGs+DQMLMTqn9Ohf4JkEqpprHE
HH2pztVeEq93RipXJcQG47sv4EzftvMhes/pPm8DfqVawMSeUZY4N3/DjiQchJSwU1iavzreFcbz
WVn2w9LO8seinRZSdKj7Mvs7QhABJvDJ6BYSLGPs7C1rZefB/vd9N8jdvcNVMY2wknc/ZiA8wr5D
kUOHMNBDVTA2W4RjYavwKNctupjW5+C6+D9RVOzEhmJAddK398/Jpl+pMoryEsGl76h4AwehDbiU
OjlDHFiJr30AFrfR2zGJjI0Mo1ULSCXJc2aslikHhtHYEeqYbUOe13PyShiWuO2DyN95HFQAusum
971oGWSUJqpu0JJXy5Ir0fSPs+ksyrxomODzzpuEHYGwJmpprIO0v+O4baCwqMceZ56v2Kds/12U
WwcyslIl/c8PL30UaGPZyCSYeHLde0JF0Tq7GLmVtw/R/z5VQc29S8o3qxreYMPajb3sVIv20hDZ
H+z/zcpMO0bnNHoXn3SN5wk9oWVL2XYPZ2DQb8bP3DCO2N/VEL5ocvXzDRcTDRo6v3pOjIHGJPNL
xjaflMvkzISah9iuDcc6zNvk1SQAaPJ82eXPxAOB1gJ6fZAE7tiYKaRRFCirdo2zhGDsibycBIWt
HUEosoQ51QgoweWySBwoEhgqDT7i/edCT2jpUBlWnaD6fOVqjWjgz0CqZA8iuzAnj9xnGZeviBFr
ir8/TiDrPqW9XPg/b1RuAt+t2J9TMGWAdA2vs77RnNabkVCH1at/t9cuzPv53SdZ8QNjLU0jZXmn
iB1FCsC0Z8yg9B2lGBV2eLlFTLAfjj6RqPxGbWnQ5UAYJqW4roS8q9s5LLPXKApyzdbuSvo256My
BxKCBygepiSLrzR5NPNBIiVtFbMATxiIJVee+Vhg6z5maKluXJKjj9cOY9L4nFO9ZFIMq1jXO5CT
V7pPUuMPiHLESLmvak0rp/fU/TgByodh10AXYio1LMOGn/3VLWB3IuM2L6FtwjLSou0bIyDXyTYs
ty6K+uocyKjlO1mbToCcZqvaoqievCsZoIakJR6N3HsCSsSzs82gMJ06YPaXEVWDjJ6mo0lfQ/cl
TNX+lXizn2oF+52SfNfRQztxaDCWRWBvr80aUtxOQBKsd7n6+0bVIYd2Zl0KMHR6srDBRaFphCIy
YOhY2YZiIZweIvgFAHDuhI1NKP5M7PJWu05ueUswL8l83DUQiqa7Br2q2yYgCMSRNfJaT66JlUar
CNOs5jx4nHZf6m3OEzOyvJxf3NTVJi+dmTbcKczOSDf322HMvKs/tiYCU3Eb1wuNbTrJpUVSpWNx
IRk/EOE6TK0fWhMW+R2eLlun8IKXXH05O/4Tzs+ZuEvAQ92wi+k3u7L28z/vhnyTs4pw4Lr/qeBd
UtE74kBOm5Eks54C4fr/g/HttaVwHF+17n9wH5IfefgJn9SAaO5g1JUzf70eGbPxaOnOOr1d6GcY
P/zHrKgO5h47m4rSG5k4TEw+6Dzavnr3BAz0e1VLzLeDsqLeHeEILqQ3ciyn/Vv1soKZClApiULU
88aduX+hDw+q6YFW1UjHNJjvx1LelqHGKr3ai2tdgn7SQ0Gctx3L7Ozyot2mEG8TLWK0/VffASnC
OGA00tPsFNalsXeY4A2v+MHSKrxnehCR1fcLa1fxRistcnlq+RfmxyI/w2lICFwCNb3pQNIqv2IB
V6ciNR1wT+uU0yLDkGX7agxk/+IvDziL1ZQGUOujrcp57HThjKTCJIRg4Uwg4FW8e8jRSKW6XRKk
3raDSQF+ogfY2rip2b0zCtX0kqiURBwBICf5peoJw6FOiQCIC6e1CI6sDy0dOL3qDdM+STbg1FDG
bwL+o+qev1F+OfN2mwA0R/OG5SwPBJn4okWg8gMcDZLSg5OZKzBMI49d68cAAlpItW5EpSf/3Tpl
LX0D/4XtJ6A0/ccgBZaT05r+2vVIcWsGeOu48VHjo9Pl3nWhXpaOqeRCAb/KNT4zIxXt56ibtJ1x
F2YPqQu4KpjFrLowpzLrIiIa7bkuoCVnHR0DTZDmz1LIB7Ro8C7nzv0Nw0eyqIIAZshY1FhWp8yY
dog9N8p4rUg45bSk7rGVwx28MNcXbAYchdv5rdx32xwej94I4iSc0BO2dxbJx7yO8yrBkM51HwMm
MOdK0ySW8d6Cy/nTVi3DkZav+t2YYn8cUofMfFLhnQF8mdaen9ZCKVzmZuI6olF+dPPb20brO+LZ
WvyaLjfmSQXVd1oZSJNE7EItQ04uIwqXmKWX/RoE++smhcmh+peXW8O3ki6eu7bW+aV4QsvJ68Yb
2Sd8wtouOoMP2k62+6lJYTKXtT5b9fbZLmoDDYpOtnK1iiGxuyoSw4xUQ4RdRz6UcDJIh/n5HePX
+2v8gqbbaGfLGbfHYIkJZytpeB5+9RvODJsutxqz407JJCbKOyGyTz6YiTi4V3lmn56zNaOryVFd
zKEs2OyQ2Btpf3NyRr0VrxVhpNi9GnNpxoC9xLzD/ETpV9XT21Bt3mnY7in6c9tehHbL2Ix+QRAP
gnSJ5IZ/RLoi221OE9FMsAN9xRellQpZ23rT1TXGh+8EqhtQVgxLDROU4a2eRx0zczqb3abLgWIy
l487be6BELu+HkF2icHRRL5/9ggOfPqfVFgpJ1wqdJpjinvebcFOuoB0s66A50UJj/YanbYKQ1Jb
eNZpU+nJWjQsGzRxZ1hzsA57EVBc5VGkGDEExTbc4b4BjTY5hMIFQW9W0drM8uRtRTEnODfdLVEq
U/4ZlEy4eoEvg9+YZrEd0/s6g/NQGYhpzclnDHjew9PPbWoRzViBM5OjL463IwEmVwAaGZ57FSC5
Ub/Kt/NTyn3EvfiJ77wohxLRX7pDRgnuuA+h7d/So1vZOrWHoQYKHvd5sNac/RGz7wn4tNqSco7J
PcXzs4RZOWmCTewzOhX+gz5X3878Qjt+hIb+4juTO3mKUAWUpfY2Z909RqQJf81T4Zvr1Pj+43Fb
xx1PKM0QOYEMYNY7QpV/frk3rxw/1dcTIJWJOLl7o4k8nHs5d5vvTgCXnIXKFTBf+emytpnTebDR
QuCGjcVyzH9618QJIgskQjyVT1kfbtp8zviwDxGKMXSvpq3+ga+W0d5YRlxw3RfkQPOoPLKCxpW9
J/4wu89QDAcAmVUXtz9qxERSbUq0vYyrYBXon8LbSu+eipeH8Wq8/LnYrXckMB0bUNxFSUtEbZLx
ublm+DEJr8/w0hTrGWEtQw4QwCnVlObA9ixc28RnUx8S7MOaYRx/9UWkizBB5wuyeOhzQanitQvS
15emiI0klnJdbhhMF+p3n9T3esYzyFVuQCLn5K6Pa6tmxMZU5R2hmQG287WCE9FOhLoY03ash0/6
YbzT/pU/318ywb39ncF6s4prmNghAJSAM3zKg/MYEf/GhlrMuBSzQr4EVV7eHEOWPpZaW6X9LB+n
WuAmzjk/bBBkBulL08pyq4Ati4Lyr44KcpS7vk64t2+wMTm4tx61w6eqhUZUC8vpCHpn+Rx/cZ/B
Zn1t/kObEnUKn5VV1pGilY+A0JHeFDaWQuXijm3jA2FIHPjDbJv09VyUjsM3/h4Vnl44XX2olPmT
zNXi4glCSWCvAgluGCriBPc6jx2CXVEnd0R1x6B6l7ZbUa1Os8tWlm1krlVibtqicGpf03iou9Ev
gs36NaPOcPIvrGJewCDNysJ6178CV6aBvqV5X5JGow7AJ8QuUw67IYL/Z84xCdTGsi4SfW6ylHhN
lrSgLhC2htribUmvfrujLwmrNel+sOxNms+dqpHeYi2awQJuWa5lEYWh5myJq0pmmFyQORZHiAmn
6c2Nl9FAfDK9HKKzuThFHXzuNLqDGzuusVH5fxtU9WpZmMXidtB4Fq1joO+/XWF242btiruBqPA4
yjOf30ZKR1gII1LwW2uC8Hryqk/ncp8nIhRXNBMZAuYteA42Jc7CSfRBPZl6y3dICUvfw0rTeVHr
6fDQCCYb74QQDoMLlrcpwhasCx5eOP/ZUVNcsRTj4SkpSVU1h/4Mkdx0ZKUD49178LTGwc9wvUnZ
Ur97MWoKB3D/lrsCbsEuSfk4U/5FE5VD505Z0hQ89vpqZqMibRgucgXvpuYlygt7r8CEQ1OllcUu
XG2whQSIjBaY3891uJHqaaksA9PzwK1jPoAGUpmGhy1rj3bOWyDNxlGZkCEospMJhXfmx9D6mJGs
9+1i7edL6r263oRSsXCEUxFh9WIXqpdXHYY76IM9sBd3cgw4fbwvN9N2MKu/xB+CXw9DcZraJVNK
CHvcNMFub4Ypq1Hx53oXCqI/9/UNVkPBZM8V2lWWfhV+dutW4hp5Liu0CQQEJuxMCeeZSL8/u/NS
9ZItHWt86PLIEFJuKa7fSpdGBbKxtn0f0PGJVvXSN5jvvaA7gj0wZz3XDAaYQQZalZvkWCHHoJzr
rKhhaHgVJCFLisePtmKEm89Szfh9zIwaITIoJcX4z2cbSk4I05ZiK0+THMvSkykUDHwJrrMBvr24
d0eQP8ZH2hvCoi3e2WWd4N7VGaYhm3LVWpXi2dDZzk+p97Qb3Ejm9pQ0T7dWmZAB56wtHOzSslQt
eLM3PGvx9Fshna+3bvXsS63WRVYzvSsM8a3UxvACg1CM1Z79G52IlvIgE4w96Dve/51M1nrS/ssc
Yq2xJ0++xTINC5dGD7W0kWf595b8WjdjA5/WmyQhfEwvaa5oTvRmLGkX4R4RA5yHtY1qcRMLHHOw
zAg2/72heqSTCaoCiyzAsjaegKV2yZ1WDSWUGcYJrNFfrC1dmHlYEKsTqdsDsMiakkA7aaqKGCSR
f3AWkY3ZCoE+KUzYb/GHuJFj6r1L+V2/m7IjKPexkugt86b2rusID3YLM5x4HIUFqJw1EK0Dje2V
fWw6ayqJf3aawEC77nYSXDXVoD6Xo3PeetBS7dxyQwEQpE+9N1lgb5OcYXlZ7FOM+up5Xv3GeJwN
RaD8LQYIvv704xYX4rs2p9W0rwbaZF0BrPdyJqLoBm/m363lQPPofs1FsoMgMQrqlmJGa+6BrEkn
FLgaxtFcDrVUQNrBdhOOWCzSzBJ6MvpJ38sk6R2L7HxPIp9pjoK3vkNi7UzL5C/6xL/Ub8l6jIdg
AU4Xjk5aJi2HuNUou6dRX+6A91t4ZXyPe3LLj5Sxx1mllsTJlEnu6IhHKsaUpHj4E+rg+0EUpujm
l9k3BzuWToYWYpiRDklWHy61rZ20wU99TPSDzgK668cpfFynJ7bl1tHZ3Nvb6xEX0VEVoW561vkY
qH1LkyP9+mZ8YUuj7VLJHI0/4RtvnpDpisLoG0gPxUbkU0IEIR29r4XPmVCQ4DthmJtv7QD7dBVG
GT3ECbcLu2+GernjxY4surluGk882u3EwCbuQ8SPoiJxRRfYdqaHriwvfbZaYu10ti271FVGx+FI
KL9uoBWgC9wwPfx9FKT9FZHUNSjTuEk1SjHhjcrP77oaW5Mj87WLQ0h2wzu1Nf/KSo8j5g4ugHIW
cJeRYpKkQdEa6yC49ELSWQAuwxQaLscvxpGu9ydgXWy/1AE21dmfWMDHJyE3bg7MjG/AYtIAJtoP
uYaZY2BHcmQrQ5DXxB2CtkVsUM0PoKt/3VSgy8hQAl/xA5Pl2RYlu9vteRFAO+BpWffHDzAtpHHW
ejgoOQYNcBuM9fsi28PSohEC5Ir+QEHZ7mWo3sWA/J4X6PiHPtFlIsUYK0/HNly3beDustyqw0Bb
Z0VeZWnm7RkJtkGXydZYXAkhTws3RRKFWgWRThPBXMGpEjdxmSSZiqTReo6HqqikGSr+lzgtJJp0
nPXrGUmOhYrlw1gjCFqMYnXBOR4dXaJPaZ9wLj9cmGNrHFH3MRr4CQXNn44ASWDmZDUc0byPeaGC
IlAESs85v3/5Am+0F0IE1/qoUBqL0vZFyANC4PiVmF15qZ8PK72L6ldT4Wa+jpHtN4Y+8W1IrHPi
K8k6bfA68GXBeD0RWyGO/LeI4Q+cNyjM7kFTPP7PwG7Wr320wERQ0WPDNkIxDX40Ku1G9cydvTq7
8jjx6WAvd7MZShTrdHGnVe77jnQZgvCUiUmMao0xTNEE4r7dcvKJaqzSFsoq6A8CEx6YR3jrPdTw
LKdUaUH0Plm8FO6FcD2XjNzUX4eqhMl/M3Ex6qKl7i/oGEZh8Qhi76x+2xIoIQHYLTS/WPWMmPeq
5AxC1TaqxzW93yUrlMTTpOuPMiTuZvx6osIt++u3BGerOY7SxlsYOnl3qpcLCQSbxnIsEr3w7veE
weC8PQdLmlKDIGDtR9FdxGJd3Tkn8RTXlLJPMGJPHXdQAV4I6M8bxBAWIuObKEYrrKknzImclFHP
vSVeSWRRvoY84IyFMgtHrj2J8TaPB6cmjbDz57t3+DA8hu7KbnKoj1eNbR9Qs+TkuIhoJua1Ab1V
TYf4QqrbujVnA/zJMlgEzim75Ydk9bl/yA30h+Sxcpw3WVBSfdp2kog2IeWZwWoOJ1myElqmfkVB
U7liHW4MITDFUHd3eHLK/dXGfvzMmRN8LLvs0vCaamPEckYTQksvg2fqVlfW2kLKKVKElhymzjkI
kNeoaxPXSzQgGKHGY2GiKyr7oLmVAvnMGQ46CtZPxSTwU8hhzUlZutDMoxCKhaET+7Wb2WqxflHs
LMHUugkahAg2mgME/A1G/GoHDM63R6voWShZex+0i+UYGgKRiimychXFsX9gHdk39Gdo8dIYQ39S
Qez5tpyOVzGBZ7xaeARkgxLvJhCEdrabsCbyADWaKoYr4VUawYlHQQANh8dwXIUNBZ/c1vLj/OkP
W8p06EVnLKV5o4EpLR+1hDGBvJMwGXTqeYrqHw7Z7h5qYcU+Oub4bkE16xCiRdyv9bjOv9DcQxV/
x3255dNa43ZdUw9oWcdISb2qvexLalv0VMRAbIsqTI7H5JcIT/WSyV2WaIcZ1yZiq3A39+CTDetq
BLLvHJW+ee2nLpN62W7TRuZVvK43SRC6Jvjl9NS1II1keKMtADrH48p4tN63DT+PK4pXspQXv2Vv
E2uZ/h/AwypnJxWUDOvHUz+apdacAy02Z7H34kyEYUjT2jOJdgXcy0XFbVA4lOeD3gU58GoAZQSX
4vwOQosXWFlk7nKmofOzuJYqxHLgtfOf8GpwZ22b95mqY4o1Zj51qDMOTcnnQgr8QK1+yBsXrFRy
KixOwNsGJTOE6knZZwim4glI4jRMaFE2iQYNIWooJQx0KzWHGv6lbKUzxn/4HRVWHKg8M+nbemnE
BdxQiX9/Fq15tOIWdh49ufQmgMYBA+01L13jIMLMxmYkvcMZb1PJnUz9FNjRXT5+BSRUuY8JuIf/
7N6FNHCLNq9VqnUIjfNRe8/ZhF/yGj1Xwur30wjbn4F9oN4CFLWklEm4KNC0k36SIwXwwxegRoK8
Rjfoj9UOvm0Xp8rycOh9JzmtXBs4wUau+ygMkTyp1HKw7ILQ6eFLJtjLEoQsPreurL/HAkpnxIax
5Po6P2ka6v8Ivc6I8rH5jCbLQhkMyJJ3OO76PVA6mKi5Y8X2/QRvN4ALP4oL9DKQ/ulvSvHet5pe
mMFDeJ5aYznuuiSv3xhEtnT4/kYlZ/o1YD4jRB7Ba4YcHDh2hMVs/6iZvX3F+XpK3ans6M83BTfc
hOsqhGe5uxyRU/yFR6EBz2MXru5GNCLX6N6MD/Y8hLPqHVrKuVL9rvDT1ItE/NDNIshsGLTL5EBX
BvKaMhTAzrJ8ragLHyTOQSPmcuGMYieV8Y58reuQdUv/Cwz1hDlC7jcIFRHSvXG+KJ6XQqcvReZ/
ih8sjOpiwfkF7rmkzQM02e5GnQ5E3bzdd0JyIT7/0LIL4qYsfvLMDwXSS4UCmngbbnoD1VjrMYyD
+zgReXX4msBXTeocgzBFcs2OoJX8UOyRLLJV5RijA6O52BUTS+sN0wQp/IM2VvwmckkkHzevNbK2
ZnGvLv01urBRE44fc9MOz1lqGLnqlCxCfAH3Js6EJ5wFmg7oh/5m7S3MfTACojUcl0RN2K8flN7r
AR8P5oThB7nOsApBkCN9VFBMarJ66Iwj3uQV/IXILWkjZSFtHWljPRTqIQvoPZQ+e8BIpz//SPbZ
UFh34QP0bii72gOoPqbV/1lTAgQPuEY8XdMGyVsX0VoWKCiSLauSYw53m6WwC9k9i/jBQBLGqddD
KBU8xLTSuTbL0OoXU56c5mhMkTT+P3MjEHb5qFd+/vZ9Cv0o7p/w0rNRcBNI4DVcluV6eZNoXVU4
UwfytNLZCNFBGq8V01PBGTYzqEBGyEZqdf0rAj4cX0besALKgido2mcNd2SmPOKGU2FwRQH5DRyq
qzApHmLNuBFtbw8Ay3HzB6nk5EEexVpoR13Wh2ljPqoAiWDADWSC4AdHklZoFeVy+w2BvJl8NgvH
bQYezrUsBXH4zwQAvai3vG1IN/hsKN0/2PkT0HdZ0p4zXu8cMRjg86v8yEwY8U6HKQQV6TjCZ9bg
dfj0BQ3HhUaEKRGVGLOBC5iLMyzW7QZ0Ar9cBrGva1TTxTuamtjDGluiLEuxX6f/5Wfz/7mxxhXD
/HhwGObHqq5//cqEXkZnECnuOhd1h8XHhPJXV1zsBovvjGz65RwMpL2w5zltffc6AVlRIYwthd5S
gcvO8+PKnGmmNyzdzoRTZ/hLTh34iJoncF2C5YO+ToKFtSdaZhjrdStVUG1ozuEoIVOSX0GhPPva
Lli6Gt1IX8dvh9BI6da737XHYTmHaRxhcXoFO/zh4fl1C6tqi/8esFZJzqEyLGtG/4Kws8OhdCK6
+JUSlC0IonMbPL0BzrROf4eFuKmRJoheeaVlPWLZMaswP8H2e73KIf+itPP4bqwYYQP73NMMy+K5
AbOh0tx49fMgAO3s7j0rIovVRDre7A/KAbwhX9NNODD8QiCQSEkeI62CZOy+4tgCxBvFBvPslDNt
/s/R1vAQmncKeu7GDeP3kva9aMbeNXV7Sl9OyfEFtfJ66VnQ0hfu2x6MQa/+h0bOnx2hWREYe11g
aEnrbKv/3iEbbMsgg+T2tc3BJSidNwIXxIf0CRGi3UQQVpkvVL6HR9YuxIQEk1XoJyFx36xTObWc
X4EfJ5poC08DZ2dSmYNkPKWs8kXIiZDmL2om9FM55DVzJiDedMAWmgqxM+lkGaRADvJs7xG291g7
XZBgkMVBsM85mwjkSeQqi962+KhhlWTfvJuCJ8ltwcHZTNAp7Q2wl24J3CB2kppz6CF89jZg3VF+
TWU1Zy8+qHVr2W5Zm6Yi687IZJHM0m5K3CEMGak+ifIufTloSBQPOC2rcMH+D32kt9XVMiEKNPt/
6BqQS1YNt+fdgXgqSeKPzDuSyez47cCYJugvaG27Ykt1BSN3e5LzVK0+Udt6IXZ2ip5tuHlBjzt3
wKWT/fQub1MWH3vQQqyeHW/tFSwqM6DpSRO0gZFKxsfDxrUSfILUyF6Vw2dZUUfj1okrjyF1edSX
bUheb9EKENMoks/v5L783w3qNkShir8TkSlRVvWceAi6b5hneKpP0jzcivDUUoHyyhCwnwhTvzLE
X/grR45THdsfXxZ7mPnup0C0462zL7GOLnI4Wj3N7I8gJfW8cCKYdaV+CGPL0Lz1EbCoKh0DZTWW
lGYkigLy6X0kUgQkB/K2ERKv80bgfb8zup099t7W108qSfVYvb8G1u9YUHQQI2fxh1iqsZjvR+JH
uoGefv5zlpAH6qd/yJBupmIq05VNNBOM4+HrS9+5Fb92G3sFDZZajCh3VRR7ZH0ojZb2gQP/bST1
ITi1qLdgGvGtSGBSfNTQjYc7KotRH6Ml0yx5UY0givfzJJrfeB4YxFMHMcJayZK3eC9cO4kUoLKS
CUfb4HFYCNqs5Zs66uyGMNE5o6R1dl0Ent33Yq+HqF+6Tm/UXHM2EJDgoxihCzd9xVQo/c8U7MjC
oY0jBjy0pakzXr+D0FRt2077AJPWkxvP+VczQdu/9d97VdnDc8dLOF3OAaR2ORsb2tq9j2VPse42
+rF4U1yXMNpuCOYiMCvWShfnifode3+d6zqFX1MyUVCG95W08oOQifevMvJyzpmdRVw9x9bYakGh
C0DKTNtWsPkpINbq/9xGYAPk+Xv76bJZdaLCf4Cxzeya0ky2sga6nlA4JuYSwWuDPDSFnAtcA8zC
xV8Uy5H619IgOt4h5Qly2PjygoSnPTAM/yUiairrCoHMFegio1Hn4Py6tag+8gUKbXBw8VlUxQYc
UfpBw97a2ciiBM++Cj1i5ppTcJXu+GUszbIrsTTjEqTCBmN9kOwFI0S8mGIuPHah/WaedC9IMWtX
x2bGarpL2suJl9g6YYWlk1qBGlaf9nL8g8hGt5q9SXC+3kgq95b8QW7bZvNfQQQCr8AWzkOm5tv/
nC/zQUcMyN+IpKJIPKopdGs1Cm9iUb07i808AQghrxQKXBUu8o28dhnFdtaIAwDT4BTvexmIaBsN
TJPpLHYK3tdWvMLLPuGFFI8af3BBKdI1ByOewrpaSngoLVhsrRVSZ5ucDY5hqeOOWKX398ThjoeJ
JStMfsIl5+CqpJ3OyS5O7QxgXxPPeEE0wUc0fcAJYZZ2y8L1PlaH1jmUabY9Xzyq1JZxQkc5Naih
TYx+kPdMjtXewTCmePPp4eKJTIBpZ38pBPpYWCUerA1nnMx5Kp/7RzDX8Kg4VgReaGHmcCCecYS4
Cly/APxyjk/69xwrK/qcx69vWVerPbhKD9hg5Xb5jh1tdquFVa7eW0TSTut1lCoQjVKqExf3gpCv
R5B5cqsnC3gsCQgzu1Mou6ACznHR9NiUCmIwOanfvC+QsQZ02LRxKkNAHCecTqKyYUZGfPOwlt2/
2Msl+hsE1SJe+A7wNBXx5Baq/tVoejyTOB89JQommNnkx5Wys3i3CYAoQf5h/guPUPiXzabcZKKR
6Zijewx2TZTzEPeJKkEibGFph8K35ZjDINWRZfWpkFbrAO9Y7EJ6pluCqavH0mx95OpSj14PVGXy
lzCbUnZfLvWjAhj/6SkV9+Jusn0ERbR8CIlufHI/kNgiEJTf5FPbD5hP9Qy3IQQ4sCMxrFz281Zw
liF0RD33MZwr4wVauLguZ/6OZ9aG4UGb6CDTMJQzGXe+Wtz6nI4fZkYuFc+6jq+F6iEJqMQpU/K8
Jpx7t6FsircqiTLWT/abX6SbvjbcEz9M/RBtyMhGc1HgKwbkNFnWKOLA/WVzijOQwR1it7mQHrKm
d6Hum+OK7686P7Aq86uGMFVpXq4kbekC8QI6HjvYCqVyC3JjbSZnNEdAqHvCtZzsYVLZzOZHRZjo
KM6hDnLoPbnf5gTS/VfWeXNk3Trxy284wkKV38RGuyejB7vAi/W3ptkdk9ht8wN1zrQIbuB6ZjhR
9RdxPfkT35sKFystGr7fJqNlwDKwRxXoY4TVT4WvRSug3a1878msxf6ENPktCqMGfbl+aQzvBFTK
hoTPO0MvPcPiqAuZtEaaFfKGpe+ZKkZmKYNaU2cPPhD7kp1tn05lDf1oOhCYTiZ/auH1GSBeMxFM
V+NwsDTNlidkJgB2qc4uBincEvwYRMpBdQIo+koSguuWZJAya0YiHD1ZzpjyxChwJ1VytbyJUJ77
pfeaJzdWg705lsKUSk6SHo3TK2r99LKoSLU4PyDzU5VmfpyrN6CnqFa4/taedpxwpwjUeYwy3ui0
798Hatm2BPrHecddG+xAPkci16W3U/GtwtXPmSF9f8bZEDwGGcduoFcGkqO2x6AjBNMA2Xs6UIDu
6zbCxN2XkkA6QYBUc6TDV2pra/nbx5eWQaTEpOauETg/YNHIPKyj/eeLBOWzOY4580QI17CTf3Fg
cOm/gB0l8JqTmZ42W6pNDCR1bcjv/piKHa0lOExVnI79O2J2hDUwukWK5KTTZ4WJrloitIEKjtoB
K9cKtsu6IjiqARtUyQuM+Q8VDrxXL/pN4ep/JcY5JuoZmZ/SAcG/OmnOHkT9mJ3zswcQDGTU+Cnx
vb/rWcRO1Mt1SpFGtYEidFNGiPXMfZhlgtCqGk44Y7FouqjNGzlNP2nNHk4tsjnneNJZPWYeXMgQ
0f5cbWhrJThRAdscpBmMcGPGhUwLPbRrWS1usswk5rj0ihj8VXzl/qclBtvUYP1ynC0uHkiB68F5
6NH3Y8yDUYR6m6LrHjs/8GhLYSEysvEcBaVrjB+2Pcsmwzm7QaDHYCDvohkRaIQ3pFA/BXLFGHva
tBIomeoogRsFLOZ3RCk5T1ldZYpC67crvBr2iR3RkWaamBxugN4Qac1U3VAmcIME7R/emZIl7ixO
p4lUgjnn7W5l8xnNbkr/m/Zkybod7A+SAtZlv4rD7vLCfoeilZIEEk+WyTRDtcyRtBPP8FGaGWz7
XFD8T+NFwkme1KiudmwMcAbS67IZhPKXq0WhpeMMBupykgYKbZXeRAQModuMQK81zZITymqEQAgc
8tvp8Sog5HE5LediM7ZHBoSnDpp8DMk5C9kyH5WpTOg6pBxrRJNrDtQlWiJ9hNP1JXzdG/yTS0QH
YD3NbnHIK0lf5CYNqKj+d1tpkuwXmO7xys8Ln3zmBB/CIZ4fqp9bXjyNLjzigon9jx7s8MIMqUZY
0W+R81yxKG00tj2yFG1shrCJjipHO36B2aoAuWU7xVcILlTJUuruvb9SVF2FE3BSe7D50TMbqSQf
cfegkN/YMDrkJOH0ChkMlPZuNwy09lM4IgJON+y5zWswf2DDylPrShqOhxNOmJMzRPVkoZ5+CBt0
8qSNCn4jcFWadeQYdqAjxcdwRvlWpow0FWPLXGKzVNpidRVTGUy9eNmxSiPr5wTcgLL3y3FiqCU+
ThNcpkQPBmLlhL1KwIgwiigT9VUCD9+Cfw2lxEp5bkBSVzwleMBDkLx0ac9CWuqXBW1vFooLytPd
PYdJPsFBqqUtc3cCfDY5nWI94w0KGkCPMNI0J7ryAlsg4ZPpioq8V5hNOEEbfl6IRUvd3twVLX3U
uDDSYk7DXhgjrfoUgylxv+ZEfSc8kHLNHnIF+XkR7E1QyOu3AwMJ9cIZNVE4ZEDXSnwPni/NFj/3
mmKBZMfuX6R8Yo78qH/nqgFe8Maro+4WdFecM4ZPt0SLfiQMmq8nlFVOuq/6B+GJ02LZcP0G2rEp
dGNox0F+9FZ7wZ9ATGc+l/5jSCwDRocAuqnHqxTD6yavnPPjXf3V0du270k7w20YUrlvgTsBP6qM
juDPi/RZHNIjhFMzO68leaLb7QvLY+ezr+XGsfM2p8xivjCkD4GgAiEs+rCv1MQzC0aFxDCBD/qO
5ansQ0G5i2krUhVWTexMjeB2lQXN+x3J2xt5hwMswEVBOu9Iz9P8F0tCIoCwXujZdtjYG9cl8P/d
+OaMcLy9pApHLfSu2UBttiVbi7b8Ebk3eEjPclq49rs4kRBjaiv5w1yEEQIhgmuluFu9tjhd4G80
FOTEgU/+GgL4lnhmJ6MeyeabxcunjlNuAXvcfJx8LyeKmESoKUJ0r3SQogZg0DsUZFQO32bviH5I
i2pePgMv4GAszZZRqYOTH0dn58zNxJoYWvYm+hwYtBav0f6nWxX3QcNQo6HImpPU5yvlvAGXGXXP
dlcqg1Zp914NPkY5P3zl52YuqIg1XjRgD0BxROn9QCAJyW/qUez9l6/STygGgPaksqR1ItyG2liA
yjWQF9LztNPPLglRQjpAokCTeCb4SaQurrUIR/7rA8+4lakL6jJ2ddtzfSoiP4d/PErqRSpIpdtV
xRRDIaOr4mEu+DseqOA/hFqf2H9+9wnvrfOpnxDjMx1CJaI6ZReALvW0CnmqwKhjalqWJM1hf0OH
Fdf8JETp3/UmDWadziUfF8A/0IorVHua29wiDZdqX6Vw4fxZrQLJQFSE6HBDWyC2B/oRlAYecYaD
+QYO/PeJU4qv93rJL35s4j2hhrZqeYNlHarETTZlMWn3j2/2dlOHt4FrBS0YjQl9YuMHo1HPlaPI
I5Yd7uOI29g1vDk4j3T0cjiwTlBUENl2M+2oiYu7WJL8USaSlyidApoVoKQ/sDLSzSX9o8+Ali52
FVb51TC40Z0AU9IBJLe+4gVHdRWKQwcNYgWlveEp1aqnpSvyJbsIJS+/yob9qwSjX7/WxMo1itn+
Vc5IofCJwjTywe0acGnbLKPXAkVJoTqfqaXA1h0j9g+HgjvWVuO+hAeVG73SDAi9pJA3vEc6Cd4q
AZSbTJCbFVd9Y9nj+56lxYmG3FIk/tDy6AMSYkGcRCt3kAtvWP2whQZaMDqqi+DcJlMkgfI2U3F1
dBvZBfAXudlc8awXDQK6v4N8yNTH5GmP9ZwfcWM5+B/iKFKnckioVDfIl06FLzDlpDKvmC3A9e/u
xJxQvfelwTii/UmdFEbdXidxxXj/1p7SDJ597ULQVDcHltsTzgs7QXmtZYqWsgNzIgCUCEEMm7lp
J7nrKCyib3NZzIE1auLtcp2ALn4vXdiMel8cB1P3dARL2YXc9C+yabhanK9QFlAu14hly/gIwYVB
hJhhfQxLhOQirm3I5FwxeVaggz9C45cNkM/D8lSHTAaMQLtvSpeVbT1Cd50hV/ok7oSYy5TzVJWK
ROKQ+oHavkpQQX9s02nh561vwPU4Z7RhOo2ryXA04R9dwJlfsSGMNXqQg3u5T4M27XsOkD0Hv6VU
xCvJuRgzNNXUeLGQg5GylQ2sz6VQLmNxXEXV6EzAlBGx9aTGU8EM2NQh1SL+qUcXk0x4sEuhSZ0f
j/Qqi7s65IlX5m/nFSY/Jh9oS3DGLjr/16UNjxoMyAdyzIJ8zTC3ELid+u3Iyc41Jnrg3NqSLxVs
Aof9458iwkxawIuPCqJFixLnt83f/SOPbvjy4RYMaSNwW2tY7xkTLjR1DxQ4KaDLD/om1LykapzY
GnNV3eg3hOQlDe0w5HRGuYNcyqOZRNtwUOj6PGTDzQ8m1J4p6inoynxfdb69FKU5DzfUkrNOox5f
DlvpJviQ56EvzlBIVbweYlEe/PVs3xlbpIfPKVxT90YaDcrP9OmLVpe5fL5oIkFrXMHQtipzYo4n
KItZnn730UNbxY4lmAXVeVyjtKLEhQmqnSETxjUstb0Jb4I2+b+Kb3DitQnFUgJfu9lIKC8/ZsuE
qBKhyxy5RsUvxw9yiZdU0bpnjWFwQHmUt3HlhNQUVrQphJRUpyi8Ie2hMuaQqqks/RdmiCegBVYh
+bls7cEb3hA4LCoVXLITtjvBWmcbZ/NcQ33kupMBd3YQiyzaQIwyB4fbQLfhl94z6CeKvgahwaKe
a1RHxnDOwDw322F0CYD3pDtp4AFDVIr8pkvSk7rCglS5Mn1Me46pdubCerYkZ+vhlKM3PIcZFcQr
mMDDiv9s19Z4O+KhM91rWn8lsxKS1Q5K1MhX6CamjSRglQPs0RncXwGloXPKQBjvjm2LdXtYdVS9
ejns6hFxDveU1vhakATj3FLBo8Np1wFiYwJ4rqo+K04sci/gz4q2rato9g9gJU/pBpF8PP5LtLNB
Bgu70382TWnaV3K3t3Rje2YQQ5N+1FOLEcor9bq1ValqgYWZiTnxz1jzjeMJqcz0z7hFh2x8QDEP
DeJ+H0fZi3kwc2igiTp6V8p+ToECa+E+sfmDtFAzxu7mkm1tGJlwMzwVMSRbJZ4DoFPZtDV1RleC
uqnuHZr4zn5tDQW33M+6AI+gR62IltKgkv3Z5fZPSKbpzNmv2h30fGukifg1EHPU4+Mab+dxCp2o
6zWh7WV3dQVa1NwwznyIXxy+dUe6IpMOx5TiVq1RPB74/RDuTjX7UTN2oGE7uIE87NiMlZ42UcXI
ZMQ6fNeUoVfxjBYA2Cb/jWBBoLwLDXjeyvYSdhH0S/piWHotEE1nEaj1OZ2hS8dZZbFQnS9ZFT7Z
NlnKz2K+aRbuC+CRUHpRONTQ1dUEh0A995caBaHeS1Wpp6BimLgouZq4dGjVrwTEcTEnXB23IMfb
Ar5R+SK/Sb2Kr/2Xl2Jxq8/SfXYkoets/yTyAO5vd0B5y/egJD9hXv+nQSklmoFTczPjsZpHFmRa
gcc5RiVgxKS5LnSU7yKRw/EBNOdcL0BpBx84mDGmHs5t8/xeH3TBHe79nSo4fPQDnw1F0KOEUbPW
Uxxk5Hmc9Q7q0IjMjJmYUzWXOf7BteOFDFxDFgbew1E+uo+WfLU5JhHDDrwzyQDNri4NQJeUAx5W
ki8Z9glHt8sAD0MGi1hKI/OXRuZhlvfB41GcBwl2rAREOca7XzgOHQNTOgm6dg1MhERubI29OuMm
4gs/WbW4+qEBozmkqkHqyk4T8udTzHFSAkMY7w0s0f9vdEtQOuDoWHQPugPlKkCzXm4PqRksyaJH
aVezzrfM+dTSvUhK66UXXBgEe7068J9+6mw52EvPt8E0s3vYvdc1QXJqQqEEYlG4f8uPTsUg03Km
W2O356JjUD5El2DqokAXZKAeXRJQCV3/pG/3taqacatABzEr7q75dbdVXV97JF11k1bSgyHEwEkm
E5w/qzCb7uQylJxgyB9GAHiZmtkqNzKWLnYpieaqnknJtPvmdIKV2zgBZWtO2117B58NGnLkVtVH
Hd+TBVJJ0/sWQnsTjukNnmZecxkMOUsGr+RBcip54LxbOmGUWrpJgpq/dLVAUQOCU5ggKg5B2N2M
FlGvaYYbWmFXZvnGHof6EJ5+XgI9yxP8XuFbTEDKD3Ras4wSDWCNkJPnEiWvrDi+DsRnLtjrTugs
PmfVdda6sKaMihJuka9T4cbfMIuSPjDgZcp15dQPh4pk38ad9Bl7ROL/XfVoZmoOYSD4AWS0k6oJ
gG/Y+iGbRPn0t9EoiRHKjTAsy3Fhy0x/V0aBaP+3Q+r0ODQhXi0WfqnvNvmmb2JjlY4Mpzsmtapa
56+9JKu9EaBOZBwZ8Fy3VMQ+jCsOutNJ+5/OMqylm4+ocuzKdsc7jS+adxpWvqI0XM7dn454Gvo9
7wgpkVUBJs/Fvxtt2/hywvtReUp8ODhAqmOE6e5jDjLJXAIToiAGOLH6yzei4EobdM4IV/fxT6tz
ufylfGz0JQ4vPQ0vcj+TPBt8ZFz4YELjvN15F94wR16gGZOf7iQ6gMxrsz4Bc5l9gEHLewlaZ+SF
xKLR9ev6C9UX8Qrj5v8iHEc2z6jBNG/yBbss5PGlwfNEOfsghzOc4/C184pKxas25Y8GdyjqLFjI
haLSvmOIVoi0Rn2Znvt5t4aSPd7b718ijyG5I2Qnp7/2pBCP9N3MFSmhw8+jyRUSd9Mo1t6y9BjX
IjclJX9jdXxkh6fVIc7v+UtfYGxnK2mCIXzgqbYFvWiqRivUMDdFgkwDfiXI7nXmCN0/1wvXGsUW
gJf1mIhzZya5+oxb5jDxonkmeUG1WZm8IxvrAlDMr58eg3L+olo49TyWcSZ3C5Vh9FNpNAUfaWV/
ofY0/jH2/mg3BvOCRQXWjzRZFjoDUn5rhIk2fR0OLLPFrjEc8KlefuhIYwWO9V7Vt2L1fm91OGly
D3GJHN9QCUm785YVkj8JTf7UbACyXH4ZbOnVE3gl+jk73Uu7k1Yi+i4ocER4PVj8WTcuezObZC5w
Zhmpb6D9a8YrZ6YiAAzhJt33kbUi21G9pivrewyJD3xoO7hw/lNoaRw/RQ6py/ejIkUJuUv594I5
2oCpey+FCWrln7q4wlkoiHu0y3n4eJxR5P3qfkWU472KvvVpZO/aVEbStVxxpsh6vzLlp3YsqJUA
CwzkBNie6iRBjVcJC9IhiNHRPL/m8EqvbRx54zQJAy1YtMtc5Jnh8C7+qDPO9cWFb+56sElkPyvD
S1K5uCKHYCck7rmU0uPHcBHak/AG7Rm4pmEUyrz7hncIUA6sgazpkjZQ5LDYa2XeDv9vOja6wtRh
TbbG6QeBZMMo9oXJyFZ+3QItAGV9KxnDL6zqG5o2YThAIpVBgfljh++f62JDi8BV6MBaRwPnZP4D
Lu4V4zqE5rJqq6OjAhbkmIOh8Y0CajO/3FSvd8ootp0lTkL9ZUMUYEJMQKTzMrnk5H5k5xDEyGGT
gOiX4R4VLvvpNs7/oE5aP52FL4MDmE3pVKomVbWBQAyOZVtI0HRNphy5X+vVyf5rgCnDfAzUc0oZ
R36r75w5B/SZaeKtNeeHJXzRq35qR5fNnFIsPvVPh655Hxvdmjv+JBtxpikK/OdYRN4pKKB+HaKi
p/VFxUs0b6x4iLygOs4x39bQLjZlTW9N6xUkPXqBLPj/hZfacZs5IJdtE8SdXKvJjkLE6mEF4vOS
dsxfa/ZMI4xIpAaDnadEPjQxPUP8UK0xcaRrmnZi6EV9XSOLgJo6zBPieqCwgITRbU0sGGVMAkpv
ijOQVRKQ46nYqofsuC3X/wxIb0DdQ3Kv3q7Z0F5+N4TNhrXE3mGIa2iuI2fEKWoG4rIfvdNF7eEz
qQ2xK9vJ+jYWigpPp0tDtt/Erd0I7wzIf3LwDq6q4q0+5V1L2BzCPhqD4STIlEVGzZOf7GDGVxhG
czBm4vYaRxPuFJGGmf2ADK+lp8vZUaEYBnMH5yJrPtBAiFPd/R0DFhd8g1m3RYyPX3QJLBt8eCpp
5SGLjMCwmU6DbFT7WbUBL+6dI/wxGxBE0CIG4G3nFEXr+xBMVb2O/OwbSsAvGB740oI1s5NZHTmo
YSJMxb1cqhBMogrUTML54ObfHJnGIX55I6jdWOejKsfmUtjqBzgZhwvJjJN2R/fYd+besJ0mmRBG
q5UWbblHhk23eWn3wWXu2jhNB5VeG9KI4roD6cJPwx08J2Y/1B0OCQ6Eey3sUCBRBInH2SodL8jG
Az4ypdEe9/yONcgKX8oourCrGPBklK1GyC2gTelPuyMjcA3hhyChUrKmDkGNYKAjVHGdvsdvSRRq
o1Z7/TcMDNg3GNjofH5u6WJDqfwfys1lhkKwYCZrWc8reNVFZ2PJh/fP1win3pyrVGxngfZ7Q+K6
y6hiHEc8gaDn0ujIsijsfbExgoRSc6H5jQuxNmWnec43diVD2SiPzkONvFwpvfrWFm2H2ghkGvTI
LUAxLCRwcOeh0Z06I0w5KqXFc7KyEES8wBAb1TgyWndhgoX3X2nenUAToLHI3N7ojM23kw+33nLr
JEL8kQT1uA/CpNs0slBGPOdTcMChRCbPPKwnBJeYzFZ8+YdaanAxPybK6/t8BC+CMW3AdNcJH4pQ
/dXa4mKEZDHNxqF8D3QpWEOqjQ/0WqlOSBXJcWOUP/FUJYc1N98pdfQN3hmK/kh4FIiK38Fi1y8Q
Zq6r3YKHvkO0XzYtbGbePwIq4hsrLiIHJehzjac5jt9q4H5Jgaq1N/Ziru2WgQJR9hPKDfhSrY/M
7TMhFd/1QIM3mIrE9gAVhfzZFrV5X+TM1BPnx9cVfbYEUK6wwo4Co7+8+3UZBeU7enRj/SqKgRBu
+pI8W4npbY5f3rQXy9stv7tXApgSfal2J8xxL9/ts/XH6VRhhZKmHO2DRChOYufUWX2z3VmoEJeX
ma+oZVLpLASSdEtBZE4H/bVaJuMs5nhoA2EOpVnouq5cgALUlnJtQFSkxueI+qf4F/SBvgEco6Uz
jbMxL7Jjjm0gX00Ar/YTuoB00HP4k5YB7NN37on9IyjH8TzUcUuFiK7sgCRBaFUi9FLIUt0j4a0b
M1kwCQkHWsSwymevEjRo6Pf1+46FLuy0AoApegOEvGLQALRUjXH7GZq87CvJuvA+iB86yaYpi61i
mGbnHb+go9d4TVn50UAAvHGzE5uh6OdX+UZnOHGLXIX8IPpfByfVjC8IErUjpVHdJgskcxF2EOkx
GVt5RGRojfcE6GG84FW9M/eTEo5UG3h4soxRB+m25TbwqziDQxF1Jf7AFM21VuGa7E9JzjPDEC4A
gwiGTs/DDqdfsZIZDy0GcNqJEiMxqSGDyIKCIg9+TD2wL70oF5nlwm94cwDqt9lUIzTVVXvZSoXn
3YJKwZRouWdHxBAkVm6pM4BuccVF2+SnkNEEY9VuwOIoypdjB1XV7anUtjAen7G45cOW+wpLnhqr
oUv75lZ6U+QI7h8GGrr/M2PrYa5p0I4gKPw21V82rdJ9he1bPIJuiVvm2mEWCxOkOkOaG7C98q/N
l9UZ79ln/z5KNRUFV/AEkpclwp6EtfSgU8jJkeHMo3GgXZVqY+D47sIXdJMPXdza5WDEbTPv7adK
VxXkwrijw8RDL1VLJW02UJnc67Nmfe2OXcY5zAdfkxQjHfFbzItw9dfWu0o+cLY8ga2tSva8PQ7J
ALUQqqFaXXKwhfIW6auiYOwztv8P3cS9YwyvvlgYh7T1TIwc1uXFk2JhnKX9zvb5i+4kmRxrWuKl
DePE5Fw6Z1HuMD+eyC6eWkUhSnEXNa25DhNvTyoQ6gPQBb0ogjcquwmuRdu2vIPNmZy/Iu1UxTAc
w+o7dHyu7heTtEES6eZSwTYcQbVeqCfnLAzkXkQFML9gZ18gOIp5J2KoA7BP6KGvpcrOX13lmea8
ofpbn6eglc6Dbts6iBEQhWOS3InOVp6urxMAYqQlqax7Fbhj0MqsV7FnmhTjjPY2eMjGBuwI/cLd
AUiD9/3V3MzTsmgu27GnlS5SQ9gNkEeiy4kvnOI3Mjkj+fsIa34tI3LOR2E3LEY8EunR4iat6t09
L3IJmxZABz6ae85YNhX2Ca4KVKhjtFC7M7xJUwHko4eMTBm+uxmfsHOLEJD7MHbUTAw50gMo1EE9
wyQ6qvkN+ztuHlKIX+RpFtkSptWJ5VKAJ/5gxAAHBa8ckSInevRMZ5Y1YjUpLTH0Ucat5LM5TuQy
WHG1CG+xwxolurK6XExtnEPfweQwxmbzN4ahxBBCutdwxIlES4SamvE/BTK83WbSHmlGRtbb22Am
X/hP6vPyAba7gVbJG9Z/lOCXIgJIzIUVrf9eS95f0bzflwS/AHNAuv0b2aYwt/mw/G/4FJBkC+2+
VHxuyJkFlOu6gMSuNx8VfFlYGOUPr0Yx25mGK5WjpOyC9K0cPjAKjIYP5k7yQLsytWaokn9w3MF0
31m/+fBJqE7avHVFeNFPOxWgGIXbZhJDjABGOFLlvJWRU7c8LA2ZfxzEmk0atV1L72UdWl3K7KV/
ycB9JrHCNsp3hsUdFR6R+CLs80Nz6P24oZpiEjYArN2gs0C8j4gI3vgvFjkgWEkBHYp88XK0d1VO
wSwJUkdc7UlgB82Te8VrKchUpPVTxoC6wNGQ320OMA0QaRKR/mUFu2BpQZgvj35WLjTgEVeUF9fX
Jf71Wh2pr+D+j/Q3B+5eurteQ7yM3SUHD/CWafQ8v5IKSjPHTU029uS0Xe4mIJCgYWUdaT2BDGS3
vSyMVFBViP2oRz9gFVs+X5asU55Mv1LL0E7V0/SYi+z2/S65W9m/Zyl1A5T42N5K8ZHkncDgsADc
k43Sj3x+VJe000w+1C11XbTUVmLHYcRgKBh+pZywL+OEqv/OkAW+TWEt/NH5rB4MmzOWsAoujfNO
0P6avR54LyKssZabYtXDvHTN1XU2e+Wg8NJ9ucxn7yZ1T0R/CGjqv43C6qQEUd4nxISwXXLYJ11l
1FgYFtHfjbN7E+5k1fWv+OkbKAIFJzUA1iJzBV4usVcxA6lrzZ3u4CyDdXmau2zlnpUjmc4ueIML
sbun8e9sspTieP5Qrx78MOyCNnjY0slXUXYcDDvh0L8Pso1k0182LB7vWb3Shxf3rAymKBl9BmSa
Ra/ZrctqaJY/ywiHjsk5lr+M6BuAluUD/xbunfOSFVpYGKHPdJ4Ujw76Et2duC8QO9Gd7P0e/y/N
M7Bmaj8oFmdFOnYz2njlhC2E6BAmgqkBFzJw5C9gmpQMk0yBXUWgaFfInO32BqgDjVcybxq+HVK8
k+IBs2legF9uw1ifVDwvxZNh/7YGsLb0XK8sA6dOxmmX2DJ7qJS5TP5TSGngJDKs+59/roFpY/1N
h1SRIoEcOAa51Eha59ETdboAaxnRECTFqHSOJg8FW5nKKVzt73B7Fxh7yPmCXflweX24w9ooy7qY
YrsK1kyyLU/9kfV+498HX8G8h4Vz23/w7TAPOlIUsD1SHZLX4RSRDpr5TEfMMNc8zrWUKloJtrds
L0Flz+vBB3Ctz1U5apentjpHLNRb6uQDwemUp5ZRVvjw3uPm8OLklHu+P/LntUTiraCPuiELUBNv
XrPDhZDamYkCaFzPFrzuAIQih74LQ6vog80PZQrNXvXcsN9cnP9tUA/yVN5mum4cMqhANWcwx5Zd
VQ3S5cpQI48mGaQ6aMWL/MUHfvgMZ9FFi0DdkDkRkcZkops7qt7z3cjg8nCQvGjgocvXaDvMxjtC
J7CsCVLlTid8Mym8wje8YdAjiFSzurLVlG7Dw1kTQm/w0fTYV7/0TKgSRMVQLrq5xnZ0RzCOPOx9
Xa0WpPnREWYwhXea89ghpgARaOaHkR4iCXvqJ6kZtlWgsUNk84/2vC6H2KSS84sFYoewJGHZEQqx
eyhtdnMFjuU+F7r8ne4NgtFrGedzHFULMfobnYVLJoUktyWN30lxrqyU4la+Yp6V/Y2GVfnF064Q
gdeDmE0eIvSAlgnPYapIOks7ybVwoHWvzaclhEulcQAd/vcx55Bd50dsVeOqRgeuvcoYo0Yyt0Ep
GXmTPrUEiHMog5xY6uOiS8FxkHmDiGtZUyXFZKGCN6HIf93ov34IcW+a4DZXIIh+foRLMGwVCba3
H25/vKht2gy6Zo5vaLJoUXjGJfcYaoHuwX2yBQb/FFV1q9y9rtYwRDl03XFSH5YDSHiZPYr0/zIJ
I7lWWASmFD+6ggrGehYOvosZwOAYvtF6QuwE9vw/vigpPIiwqbf3zPDYPHGE3Yy2MGABSb9U9WEl
1HYKbKXgZz2/naNrN6bBM27iPg21hs7c9vK8EpbLMvr2PKeSrlGizBQ9r3w8E/6pv6pv71UE5weS
cM07NmWSvgLJ07hsfvu3cE7pEj6RYJjfdduRUyA3kQ1X5oxcYckZURWqag9gxFyQn4Rm+Pj3NR3x
XuetOeV1ffMkdckZ/BS7BCUNDFABmQbl4wbEgOVXTifLuE4icYyT7viI8wAcj6A/4zn/oCa66aZ+
NuJaDWta4KjkBZ+pIAD6xEcstP98lt2fpvWMZ0c+oDwp6enYs6ctaNeWGlWhnfgRl62uItj+DVmq
rTJl45TZZCGqxfC58GtojlHLGHl2JdXIQbQwJcLsRpN9WqdkxBHBYIMWdi/hrj1lL9+IldwW8F4e
onqq2IQ/I4BtjPU9CB1rR/IEHSbww3smthAKYE6j20nzZcfqgThasxdFked6c9j8KLike2YiRQ8x
+uSxaPRU/sQOSJHFwk2MKjAM3LyYH84n1JSaDN7MobMx9/O2VD+yER/aVit4QUxYB6cm6lBoWwCy
MxEhTS5HD5qs5h8yZTxKzAz4l22Q4wtCWV6YXeGX+iyshlDpkRF9/H1wP60zwwTpKoSmPxm5/htO
bj4TeJWy1jh6AbxHLZsWnPA3snkuPIl76yiZihrn8SrqrQwzFxr6xmyeUQ6OaD+CeTgspvHbfIz9
qkdeIBngYn8QzdodecZ/o2Q2VLzPNdxBxFw4J6VnlBY2WUwVSh/75m6kzmAJyFDVnjuctLXAGaZG
coBG7vKIGoVNwY/ific2cLROPL62ukD7/N83Pq0IOfjRby3pgTDEzKY3ijlbYh8QlSLYNoxGbK4A
ymqMY2gJuGrmO4hWX8IoCpGXX7E5i9Y9Ql5f0hzQzLJ1incypxOtKQD3YTI3Ila6lradUEf13D8W
aGDvc0VcpnOZNpSE/eCB2AJ8gXDTbwWwmuf1mH7YB2equX4jbxGR2aBIIdB5G4Q/+Xf8kvHaXmJ1
w+pFdyAkxgONic/UXuGsWwLJivzSdN1wLPnHNJiQ2t+6K0Lvu3rB+ALFB0qZG6jKEa5MszIObQLy
gGmH/E2X4TX6cV/8KenX3FZ3T200imjvifnArPMP7qutRfQAUx2TKFQu1DLDmJb484i4BR7XDqvw
sG1TXeHZDj20F3mZCl5wAXZsrEMzUsafOAGlZqzIHqFTC5Rr696dvC7M/9qqw+Dh+GsHnSNEW8M+
a+GFtO0+9KnDMvSjmJ3w0PxZbKKa2dyt76PfCSFr0wWTaAj8Ehr1JuGqd2fZfXqcfx26lAIHcyJS
e5G2pAgvwwm20kvBYWTZlytKPjQ5BsOhwoqMxwHGwo+oqjiZegmBA+riGK4HJ4zpyr9UoMhUULwC
1vthGPEzI0x9sguxLa1nTAqbOzaq9Aq2D8I+umrMPaHohhZutAAEcXLJzt2PfZ9BC/Yo2vx4FcST
UsNnAfBFEd9vjbW/FxysAB8NfrMb8tSiorLuFYYpzYLzna0YFpP28iCVTFqZJwNenLT5ByKMs02o
xKq3afhAePyvnCTLGV67DStUxfMd6JxRjwbh7zraHzKmVUjy9F1Zpw7PD45BEzQyVNUTa5jpcnHW
hySuPPnQC2G9iY+MDE9k6BPgD8o+dZeX4LPhy7XVEJBxNfImbt+TRyg/D1zocJgTggtUr8UPBWvw
lvld34/U/Fn0I4ojSfsf00Pa+TGknXVo97+N6+fdZ1BgC/MDKlBTAiaIEUIEWIGaxKHYZ0sbZwoX
S4kR5eScM8WOzHcIo1LUfCJwSlxQ6ZBKCfcP17vKS0szJFzHFyNbsEfKme4QEGnJ6bcBjOYKmZRL
8/CwQDFbyxHtQenNpuwK57g0Dx+OX1X/b8XVkZxWcdn/PhOLUsGfc9c3OIVOs74gwG3tKrYLStCL
YxHDGToB6hW6HI/VyGRg4yheL6lG4BnZQReCGF6ND+xRiqzSlD+B8aZZfPShOgLD7fm55Fvx3+6W
JinCkM32DQ4frf8l5CWJUUpcaKUywONi1V4sQCzM4dc6okL0QcrCq6cg4x0xrFLCNPdPDqHW85n6
BYX6JPNsZ0AMpaNU6OZciY9OpLumXR7Jc4UBG+yygsj/cuL50hmrxsPUz01X5B37jBeQlpI7+uBG
PreS/IfstOgBX2xizPV1hgUUPqL7+xVI6W+yCfWfS3L5Su6W8qttKiJhJlHyO3vuy1P5Si9tz4/m
9w0leg+KPbvA+zDSX8wBj14sv5HAsi4bL8YAa60/CMvWJIPjrhZf7mFnnUj8ru2si36ef91psQRm
Ax21j09xDOWFdTSw1IrxSks0b8AvjMTjJg/eFG6q+n85+iXM8UbtYHJQHyPTVMM2L1akygkDQhFZ
s2Hp/WWKmJCprTT4ureBlBAhBDaK3YR2MYqhdpjIJl8mHJEPfJG0Rp2VUf6FHJC/LIkOaCOuP5qC
u9V4H3RZoK10fBW6gbm2k3cRzK+tP7Tq9NlwR+XGzuhGW1u+uc7V+b6GYiL1NA0RV6jLAo4UnmUU
bb+iXxxyLovc5YwzPgWqQW+mxOOPmDMK3qECJvbP2Jnq9ZmZnZUX2/RfecsOtdhm8KmNEeJNWVuR
oymzqra5Gvto9ok7jdxdVNQddmpywrtUujKkP2DDAhVn0bZgglI7s659vYCbOgVF7OfyB14AdOzO
pGVQIOlSgcba9/VldLJSyFu4oLRZi69dQQUWOIFeSY0xB6ybY0GM0GY3GWG9OF0nXTl+YH/jr9/c
isu+Co+P6mhzAPOzVmMyZNuMgDUJ17WY+b/kyv4m4JlgSxJwMC8c7OTuoPvhP1vpbKTOTGjhQAXu
MB9uItWXnxAXq2lgbPo4sOFYpv8+m9fhlAVad9UTHq3Gv1l9xy11BOGd9JRngvh+xB2C4ZuOmql7
Gzvds3PxC+9Aocl3giatcFdNoGrZwPtzr0xDS7dVUAiQ3PaSGuVmxvTTq5SUZNHmuEUjwAPFeCWz
2+slP/Z8B2c1Ole3S5u1qDQ2wjalgbVKH+H3hBjTAb9XbBYbJeKkXzDeE75socYgvcGmwK5qSdP/
S23zBkxvGexikVGgEZsV4eCciHnrGLpaesoMEcre8jSbpmuj9Z2vLyEodesjOKuGXAT/lKiPmObm
raBuZo3CEf8n3eUljasMGaNOXattdENdqqwM7UMkwfKCVVYJrx+Tzdq/8Kfuq0zYxcVQoIqmb0qA
Ld5BHDSrJnC+9KHI1Ci+BrN49jnSIWnbXgMVpCe41EYcW+bw8RFHKx7DJTdr3cRmjOS5a64lXOzH
OXCPkMpug+MmZ2NeIcCNgTyuf1p2W0pPLtLfQBmURo0DePeLzT2YwOv50AsOIzI1a5XmTTIzG4SN
2u3IL9y3qcT/VTWShW5j1QCX4mwWC1Pw2C7m+mtHGiF97+sMbdvsBWWyIxzs4oRaS+sVnR4LfyjX
OEYFbyqkB9MuzxfN9hKPKnrpg0mMi2lXmTd/y8N7W1hjdIQfJzUFQo10ZAnYPIwo2RiwNW4JtzEb
Qqcf7LNdOpzsYhoi3T3GCdJd4AhLhjqOIlFuseaAP3UeaAPtUPnWHyB2Zl/04eB+NFIq8GwwM27R
0tbh2C9wqqSYaXuqmRe95FznTTQTQMyuzTD9pKVfID1y/pvOkk6VwW5p+1QVSrhoCvlTUy5ERO5f
eiMYsuD8H2cw5mFhw7vTdxVWLCdOdRarDHRs1Wt0D/wwH3y05gw0GmT/EbfIMxPP2VwQ0O1FyV+O
9FABRPj4u+0+FQcszOYBzdUICjSY3hfa1W3a02TpVSFChMykTwerERM8CleMFPpNvtHWiUIkHsrX
H5BmAOeuGzq0YC3WYGwLkJlDS2oBLdTieGjsYY7OFBiMcyFLdWYFxUkpLcJCYIOn8IPMJdbsspcz
KUgeikFZ/AmX8/L2ug/VfobysYw5Df66pVmv9VpouD/ptdLo7kmZd3nWvOa4TiJR2QoQMlMPjfvI
1NXpWIZzcjNBO2Ir5xTTT/3t/FZKEYhjIYS+KZGKgONWOXiAxxeR7DIGzKgYjAOZpH94o2mk9JnG
q1gCArk6jv8IlP+/lgGdBCqsfnAwgn40OjqMdkwVPLVokChpdwLuluq/o6DU96fkVUJ5w0Xfaszs
zJJeB1vqJW7iEbFlT8UGYi1ZGecYd1W85HBYD416Mfc23n/89oAYquCDu7TcQ/sYFOMfTjCXAxfj
I+MFIos7voI+su14Le2XAiiHwFKfW0caJvzBbiX88ctBqJ/tT4Eg4PdWaSkQgDE49ZoLBwgHdEm9
Zct0KqY40C/CFilQnIksuRhEEB5To/l5okTlsH605C2jLIJg8s8BN4FtU8rRs08CJpTiEnzzlVFt
6nZPKND1KwMOt/aYlh5DoLS7t2cxQXUUutFtD0uO1Dd4Hk5/nuxpr7w+L/Ujh5Bo/KMMoZ1BYvRZ
33ehgXHP39gRvqN0vVCJ4acFrA97+ybM5z1gFQZwGK2ntTl1UCz6KuTrmnGDiH5LVJX/uLpauAlo
7BgvFlSk7Me0B4tnUFVP7j6vouX0N/exoXQ+GY7FbZZVG9BMg/fARyrleekuTgDcYTqdzbl+eA10
2yG9NGDC2osIQdeJBhf/L47oEASNdZFy8OK2nZ8NzEHsxiqcqaHpGpqWql7YyTrkeUsy4n6pDJvw
4exc1Chj00sPVzbHnrargjEI5tetKOMt6/Eq6PJNI9neNbXO2cpYMxzJ8W6oNhEGLvwOMpGmMmDE
RcEmuH1Pp7Uzzcu+WCSjRLBtsLeVzUAFHSptE6AHPlFPra4ToS04i8V2AeeQu9q5Ols/4y6k6Yyz
1fn6NVlzQIVIiRCBoUE+i/RLjZOH/ZpmCVO1MZG2+13NBh4KLZxJaBcG6eGKgaSr3RPpPPw90fEh
H/JWHw3SVheSWZ21nekhU6lq5b990J+VUr3xigCYg6RZaC6rV8Y2WMeCZ15ARJ5rrnzPw1dQhJAq
P5dV/agteSAJgwd33/ZTLh99hgc6TBQ70uCKeyJeQz5HYq0kGyrwbk7Fx+CrpEF7zK8YjL3wfUjK
NxQAipo3g4D94J3H4p/E5J7pgUOQpb0SARDihthoUZM8Y41HBVg9TzEv89748n6JXhqJwNMBUXKE
E2/s4ORHH3SUd96P4KxbjMZosNvE1CokNH3JjBvEtsP36B2uTmMGh99XTGiJe3mSJWzcMVPL2WOv
z8dq5NQxc7M3ArNx7alBE+6k0Yolexsf1voKM2uxKLw/RnJ3CpaG5GcjXYqs48+KQDcPT6SZ5QJi
aYkl9xtiEAZk3JDxfphYwwx2oeEu0rUEhfkxACIirufeX3yYTvVSVHElOYNz2GwCY4E/efJ5iQP5
nDExU21O2sBZJMs78EVwxB2dMUjTp6LB7nzCJYTO3jGaXifE5KTtrXKuN+CjOL3TJec05Ckm93tf
0em9BHJO0VJVIhGVj1UqVNRLei94gbe6DMlhxMElGkDo4yOGXlF82oXszULpRjPjNB8+LJTJhgcZ
zghzf/WEzcvx0zj99aZ0T7ghAA4vLMz4HNkqf7y/8DXsgcFh8pAVmwH+w0ENdVI7dRjQs2XDyV3U
QvRdYoQJQRz3ZrL9BhBGu+9XitQJpjgPy36IWeTh451hUJm94Jo0N3O7eIDRpF7Lx33rs3Nxj7Az
DzcFUt7z5nUy8n8BADbe/gRNUapURUOWSzk2IC+VVwJ2bhpD+iw/xYAWRFOVTA3bHQT8MBf/Z3y6
TfhhZjabbzXX2I1BfHHozJ82BSLVzi/2MS7NNXWdTDo6+zbx8x2RhS4RI4cNmJcGRIhe/hw3TpB3
dCsvuqeiOwzQkxJGEnv+zAIDpC4IAbFg//Iug5rH/dDnnxYqu37KulDTsWSXnpyCS5jH0uCrU/fv
jcITi0cT1HMFFyxtnxSoxyU8CxG6xRaJ2SqDhfPMKpDQs4qEgyrLHTg5/tZd1F+Lg4w/Saz8sNgb
tqpgoosLMxQNMMYWJ5RqYc7pRzNS1RYMQUIT8F3Yo6f9aoWjm4DhS87yF5TN7cf5VwkZKgo5pQXj
QiqcN2m+kFpZKJxGRGPfH7l4g0sIYk3f6FYVav55lzbZdlhOmxXflm0eQMnN1xmeLNPIMIIVoRqE
3CcAEYk14J0bWg/9pYDzWl2eI5OwwdF7AoWTwFnYvpV3c9d20m0Frtqv32oQnnR/DLtVjJ2MN026
P5xLtpJEV7n9heU2E2tL/6GKx8pKLs+LTpycllIlX/1C1nSxuaEd88PTvkdGF0awKkMTCcIERULH
yO3SUMV3LdHrrmXkwEtdisXPSlecJMEiOaZMQRhGpHWr4q3S8yg/1V8D98MLzmksy+Ri4V5Rkkdi
iYiFUg4uI56KhvZTeGNO367WkOww8Wr8eroNDa1r7mO0iNrSjfkOUSa139y0BMirTCuZYRpvNVJG
YbSaXKvu+Qv0sLesORZ2zeg1rKMpU+etMwqs8Kh80dTyGsDzn4z32A8KXQXZf+/DUHpB4By4lzkZ
d9+XZNrdHzrhR5+P5WD/nTlPnx8Q2Ob32Sdf0xpvn7x34ii5PTh0nO2TMDY/EzJYeCf7YXtYrvCs
qCpHm1DMWDCWJQjQjqYAYzBF3uLyBa1x3uMwhwzHD7e4xhHEkVTwQ0320OQmEpiJqFFTiEN5sCUu
yRdm9c+pVufdPPwSB5ruMiGEt0IGgAlUbQBUgoQQ+oyJ/SrElwVnyldyA7Zm2nVBgBboQVgtGFT9
sHziZoZt16drWW/oeZ8kRuZIXnCPpDJrLF+RdMrkP7IKGa3Z2uVuCXYbDfJgc6lVjv/anpt5dyC1
+Nvl+ro9bK/QBgPY+msheA7OYWEQNjVfOYTAh+ypoqZ7NoAO+J3Od+7Y7OJ5mBoYl6EYZapCS4WM
r/fgsRFnxE+hWX6F36WoCr/OziWVxN7QL519lVoS6bdVw+mbFNxAiS5glIVd7E4JWlUMc16xkgss
unZWPNPwA3utQ19OhsgijJCiL0EX46vEFkjNkW6iLJ4tSiJod3P916gBbgqaU0oV5quIQBPvLf0o
1bx8yrxh27YnNGrhet+GTz9nGZdKDl5dQgc3Y1tD7k8mi3sOzQpDS+AofTDV8SDbiuvg9g7+/HeX
8JZsjBHdSsDJGECBYf3d9WpSzgbFRrcu1vIkJyYkFwjvtbuaqfLkrRwYoGF2NxP9j7DGfLNj0Jqx
GREkB+GsryFnuhmcjLQv61nriek0TXc4EwsTX4292OcayvDeyiPUIt8/wCeioU1UAK9kBdM1JkbF
9nzp/fBzrcta9NbR26HUTLXXFudiV6a61oY086M862Hw7zavz2sKEgmRi4URIy3KcKBdnOhdH9kq
wNnGztQgz9dWLtmq/2axmlenjNi1bXZKNSDwXPtKHeWJLiiObkFVhe3Z1KCMbLDAfbiiYvjejd2U
nb2nwLxj6BuCe/3Ew6XgoHEii0Xb7dlNAnU8+8sWwbRmJUbWD4R6g7IUEGeRaHFKJvMJ9XWF2qxE
AdCrOVzYJShuQk6VlvmwChl02DBDtRyVE58yeFaAysMptPn8nRu3ZfMYn8aIyhmiIR9k/XJo47tL
bzrRoD01L7roBFKasfHksIz1nGPGu6ybHgKLK7hqEfgJvjSXsCVBWgwQS4i0wYlY48HzqJfNF6rW
+cRj6mquoLB0fLehQQLiXkmyFZ3aV6vIEXjW801xalhHIwSrq4i2sCqxG/lTFSnalaDcn8i7Lp+0
HmL0ylCz+ZywR9Uw3aY6gtzpZo5y5u47Vmwvb/eqXsOk9STgxquJg75zYJZfbXBiv6NrUcBz7/Ui
bzzQsiVJF6xdgcX4ACiPJ1er3V5PVAjsw9fMBEfWoO4eYAAMrqXU6pkv4rHV9utxy1CSb9aw/1hE
7RTgf94NObbFYNCaQp0By11pjJOENHSimqXm2mQS+UA8ynqeIPQ0pM3R1Gux1/9cG92Wh5IvRx0m
ptJdJLYLRCWQad+Sm3Eg7DGSy7b7QrlrnUHBNGCIpPQ6pAo0dpXlhWqTdskpZ2IRB7Qhyh5EOrfa
NASHzzlVr3qmIuiJ6PTeSnh99SY5Db3mxsGYsJ/KwC+iGnKGnqPlEGf/EXWLdTZ4SKbSZQ2mE5Um
sUv+WtWBKAxcDZ/DQSZvsmUKv3IeIsG5xtWWQmlJyQC3bylM9dpuoma8vPTgcuL+vesUz0TwJhPb
kx4gFslT21GJKCj6qeycMUa5W05aE8b88WnY6FuSX5zBWXyixh/XpebmkRYFnvyfAM7PkfjFXHzj
MyO/vdSSz4XHtpwK/2d/cPBacx4DKMdTe1xXHiZ9FOAi1dodZL8XCVyP1rGelKklDI5aYmvPpTz1
UumJ6fAV30d9d72vMN7s6gBqMgZatNlbFf3nQVLXIOQRfhrM999fdkX3RxyD7SMuQtXOHNarGT5Z
WHfoZ7+iCrQe5qgVe5LGQiXmJPlQ1deJUYfcXB9BVLtby3syZI6t8MMb3DZ/WFi+CNz7Vol1F0ts
Tn4KJyjyLSgeX8jfqg7B4b0MCCZM2taayJAwh6nRFXEIoFl9s7q8llFUVP5o9mI9Q5t53ILWOtPT
owEi8LyDZ8dqej/LnZw0R8fv9BOQBYRYd/6/YWYCBc7pyyhkQMZLxXlcpbANt0J5ZjcEu+mgkdKh
UW3TPo47oR0/yiQee4C9s2ll0KXYCKsa05zd6yVGqydf9oZ5i+4lI7QH3kVQTPDFrCC6x5h79kYd
n9Js7Wit2XIAFMenaZh266WEomU+obx4U6jkhICgzQSDv+cMUiD1J+0LejlDLdTD0AtkvonnCmTv
uDp5R00n7/B2/iW5tQdrz0aWK/jax0JPv/35tXzI8W3d5B/2c67sREeNqP5HJWGVF2js7LCIy1xf
HzU1kaD57kAsLyLafKGEkai6eOwPLFtuFg5WTwZkCADZ4xTONWNSSWH3czRwD6R8mj9CXhCKNtnq
yXUeziXBvI//PT520J04jmXqvGrKcDOn2PZpKTy/1BR4ZEdUAgq+Xa8KdJB1aKTdFq4GZkaLgZ2p
/EXxkcImiL+lMqRKAxdOBktFRskZsslUk6hAjv6wlyI0tE9TLJLBCXo+M9duokXMQES7I41wrIF4
iIUr8SuCvxDxnKtD3Zt0Eqv6fYPl+6MvrDmBjxhD+S1NrMERUEKr0xNloa6WktvpVsqRpDtfJSZB
Jqs8kOXCp5RnbWSV4Mn2Dwu8aEuaYBt1QbwJp0Xdj47P3vosETNrOHWuSFjzVOYMqcOqirBzHj3X
AmDqZ8NweKmWHGh/iwfjojN7DyyewqBKG+Z7lioJdsVmiqGlqUtUqM7zq7qa2+xm7ZEZEx4NARTM
/U6n1ZDVa66Eii/Ye4xOKCk9kV1tZd9mMiY2dz/DloJqYVfo8jCE+qwV/hNdefxlwTMKEzAbhbUa
+PjCeKnUL1z7hHdcI35s/iVigQDQXzgHSKh6NSQ4n6yKY5+eMW3Bojw33jzT/bdn0gP+D11fQyJi
EK1Y6GRZ+riSQuYw6wL8xYpIVrftCt+c7wB3nmGXITHJEWHo7yvD2x4FHnGJXvNnYjezWoydaYsg
5/OMoJpd+vLAw4yYw64yImnGCIqUbpjwqSxe46NmZc4aK5kmcRh3an55RRfv5jRgZlRlTkWWEXaw
0VqJo4hSzW7/ju5iZQjCvVTEUkfwvZdUaaduAk2OEJxfABo9uuyyUFFzThLb3SY1fuy0MG70JluS
OKNoWbl7aFchs+2AjZVLKxmrfYOV331jg13zaqcokLHyWmWsMtAXqOwc6qaQjkLhKJz3yF+x3DoG
UvfBPzcl2p46nRVoSwjnzWAtlASymbU37JvjVKpBls4vY2O5LgYFqPgj00ISoa/TkvkNoFDsigq4
Wox0d43NNmJp0bvdfetkwbIICgfeYY8xiZBZrTqvT7vUT6jF8y51pC88ETgDDQeITPZMYbAt4ooO
qiJpNDIJgRjBGr1vhunkeamJe+FOG044f8LvvQOooIfBCxAl326hw1oAeZfoAhSY3wERNH0Hamno
qBi7PW0sLJn8rLw+HleKbsCSzcIXkR+uxY6iNesPy8BQL2wED7Rc0F9b4z84UeEm9Eu3QDWSYszY
GEeFbYNHQs5lXnYqohrv/1wkkubUgnHeHgFlEg6WQxYGYuSzw85bJzPasoTIzpBrt37Wf8DhqGHP
ZPD0HoUFf2yQ9KX1bKp3u22zdR5wYdkB/xlaJuXtYEjUefNVafEUeMGwe3Orn2OSFv9Jz3+SJzxF
OJXZjhkiZhnEvPRQEFXOk0L5KVoy3ZFiKXFcunWcLtUITSSzGMQH1LaoNykPo5tTjPUl1svv8uBz
4Aqh4Z5vhwGQMrnLbbi5cTGQup832dQKb/BbxDuEFZq+OoufMeAn9HRaqQxb1ww3OMOHMpDSTf2X
b3q3aEgLUEPrVDvVK/nxlCFYuUysPBUbhTgwWggUfyffA7RWR386XuQjlRllcdk6rQ8ge3oUhPcn
OiJI0aqCZID1N+sYX9LFp3kNa9pELnRVK5cEXSqiab/IhQnvZcy5F92fNTkmMjPMchMXzF8YpmhN
oxtPfIgh0RjjvBf0CQ/5TzpqJVzS/eEtas6gwf+gsj8s+P/7sENnFwRBgyLnghSsdnaF+nfDo15f
K7h1nmmg6SCW/vHZ2GXc/J/PEVFFmwW9sCPMqhodIlL3lkjSAVq/K+Z0TeezBSaK0OeaQUCQBMhR
Qm8UIXsBATUtcOp1X2KKPB2aGmAqXxUVghVJiFRwzLJEZg5FTWzuUJXAjAq+Lr8xbxBQbQpMy4ki
Qhdy6GytUOLAg+LTlL1HjaljabJpcvds8ROcfiyQa79s8uGsPT8+t9jvvyQQH0facqeS4/usn36x
q8URQQt9CbFpNVkr6wOyjtWZxOaU5iGK0UN0cHMjDNvqIdn0p+94c3mD5rzWaOtl2uuyskvSaEpc
PslyZGWyJkQ3a2SxnaUHeSjYaIsyFYfu7TMZq7t70cWy0b3O40zHVZ0k83+mcunD0GysPz0Q2Msf
+OByzYBkh+jXD+AUJo/9jDKcNAz6NLJx4/WvWr6tLmG/JsgLQm2/8cK4SvR/D/YwvD5meRXlUdbj
WdDlsQcljbwcuE/VuXh+uebGpbefGMiqVnTI8t05DRTDlTx5c5iO8c6Mq2BimAqKE3xneKf8lxT7
ouFVwlcNUw9bOsfdc4Id1auxESaLfXaXSd3SrZ0dVBgKB1nM+pWkxbfBKfZNTXqfSgS6le0RCuHA
FIW747nWFPhd1gUkJWHH/dcveKLxjiytKwkcjb6X/KF3NRkx/Kk3Ua6V1+NFMU8QRELXzBYIouyp
9rxVYFnCLl0EaNXD8Rg8GvcemdhWZW5UvpaRmXC/l+rXFg5osqXFmJ6IY74oXeDrn5ydjyj3jnlK
BdwoTrF9qorOy42tHHvyds9ZiadyoV9f1fhigLRmVcZ7rmuQdqT/w2fMWd3O478g+vFuZ6cO/hRN
/+scSlusXCfu7ZIbN6D953Zx+ee2/4gJHdPAbk7W6rjdHSvE0I0rqogNH1JCQBazgQfFpOVOO1Uj
HrcIpqO+kjBjxNBSqjCqZqek6KCAH/ya1Km2VmfLl3kKUf66lEXSm07Yo0FR3B802b4i1XDWN0LO
L1ZGvSyxf1PTECV0KGRHfx9GkWUwxBWZT09euIzYXWyJWk9o0WrqpWrmJgHy5f/GmnNCkUifVnCV
fDPvcJefMWaqzfwV+mVMp/ESnRG6Nqd3YQIlx+DU7ZZr+ohq2sgR++2ujxwzau1+HPAQ+Pq1/bVL
XJFz5Jf6zkE4Wb75mihF656ZGSUS1mjWeIHEWU40yPcDjBK6Bvh+yb1qSpO5miKKrC6lshhWhOat
jwvZOZOnOBbY3g24bbxG0t0+oIey6zd10GLSW3SLXpGduQTl4zL+53iLK0eqbwU/NIg86If5lrbO
+L89cy0j76cS6q01YmUroNLEUfCjEoJf/agjrmmVCbbW37lBK7zVlnQrhzG6mtqZ+1paN7pzY/69
osRzVCvSsreSw8aDLFMl+1bueJLAyHgEH3YdQChjW/Kip1nQacWVlNXnaMTtUL3E9aAIILa47NbY
hhy936qq+VHo0bb8b+hF94h95quAuWXWvlgJ4ygt/L/4MRrN1M3HIyg29PMCJtidSjuyBRYT2LUh
FnjIgU7onpJP7UcxjQUrR/rzNIP/qY2PoMOPAZ36QffgiE2sudZOgxiTa4IT+74in3FIj1WHAUjH
j6TNzwr8leLutBjOdog/GGkfwlso8SyrBDZ81IC9K5fstk76S5EmVDP704kzUria3t0n9Wecmjwm
Tt4gxpQ5U2jSHFwc+LNnW0T/y8+75456DYq76eFEQ6yWHPwtT4j4jk2kSwipFXCTAu+P4YAVSaiT
pvXb6eXmCoACIQS3ojosUxb/f7IMWUwpeAOcGYVFYGydc8jB4uw88jQhn//NzeWOJt8PDfrr3rIz
aMLks0NcuSfHYRU1yClzDZ79qmFLe88GRPEhCnpNSdIjI7iQn0PnllBp0TxI2v6u+6k6gnehAGdi
9B5q3RELqNRHavsIJewWYwecKQlzvT6lhHYpGQmia4Qchj7/pEzY19xkM5IXdAtFlNJ8Z4SNAQRo
tTLIk4bEGRm/Gfg4hebMauUM6hCyIgNgdPtXMEPsqBK/sFv67P7Be+50pEpPSB7meC/mSUONI0qN
WlvKn5u8hseP/cCgx3+ktlnGakRVnatBp1cHgE0GEzETgE2z3tX8t43Uv0V7QaI0qzuIOnwaGMcl
t6PLyeiVAw3zC2E9/HdHr2Xi6rcUni/h1HSpeTJbQUzH5d1SjCaFNdMBXPMt7ite6OQpAdcqi2dL
RPYO4oUj/zEdNVAXnsGcuy3bLM62Rquu6RL+P09hMi3fafiFpVcj2+ELtn83qyxvEKqXvtFAungG
m82OZkU4xTt0RHbrHehRkb7ZyPmVQXYIzQ9P/zRZNAownACQUS2wD6USG9Md7HvyqnsQ6l4x3EO0
sedFUgis0ypiKOUDuksNBn21FvM0r5UqZifdtDN2zROKG5oz1udJW1QWrqJ8fxO7cl7YTDsBNHfz
qaBDNDil1mtK0nwLAghvn8WNTKbWs+LgaNHoO/Idqh744wtfl4EVdG4dr9Rbyw14z7QyJbLf8xDq
JNuVrQ9aWFw0dwWn7FC6qzbqCHJC0hiKAt2JeWZMWleZALOFD9CCkkwFbVgfVi4I38JR3uXpFSg9
43dYIAWqVtzgMGr+seBIy8WxbysJwQ3Lnnf4rZN5rioF0CuUCFKqrGyrUJOR71jnl0FvZKCsCDvq
uGcXXw21ftWmiwlrJaT4SvivkFGUcf4uDXXDVPJltXhLiDgMJYahzQ0c+O7LCamgpnW9ZmWwFr16
3KCUaG0g0tvkEpoM95PxZQCwpspSnpinOgk0YO/y/3Jd+ykoTTqqPZAJmB0pxZJVlBRLYDm3AzfW
btOik+/13L3KZbx9ImI1DrQ3i4ZCVIsIfz5qZIoJWai+L5WJTp469fdOjSwMU+y7xvx/l3B+ayvP
Dwo45ExY1v9z/9w9S+w2AmKzxbGBXRfnQbJHMt6IZJvTTZpoyuBOj3nCSPDO6hgGpiRp6e7Ja7Vy
3zj0vsXmxlobJmN9nZNH+5RGfJMtd6LW6CCbSOre/zbunfAp/INYq5E/rBCNDUYDPZGfnRJnIBeT
WmCtytubqpkjCPM222r4D6hUNXRQ+o4pnCUrR2OdOElg09174AUqLSJiy/AOWYdzZrO2K6W4mTfH
6ADtdALp0JdMJfL4QX14v4NTgKr0vRG1VWIb2sCAeY9Kzde2jHPOZG12P/iUWf/JZXx3ohjPuYHU
OPEb2asq5AOaHESkPPy1xC/sg0i0yY35tVkGCpTSmrESoHQ6zxnKYcGhEI1vaoy6pgBixO5mE+g1
cGG6HJOCDdZ4UKQQAfslC1Kvguuhj2zMgkepXzZp9ajtRyLHEbE4xNkxjA3VD5m5CHrOfdhCMEIc
9as/qLuOvw/aihfBKqx/QhMDkzwlh8JZIBUCeJASDp2spHMbD0Jxrzi/qen/mwQwcP0+uPGof1DD
COEugh/75FaG6qtDpItAraZmll5lfnkvfNguU+b4cJfoOtqjQqFDalfQ/rs8l4dOzAumT9cbmumc
/bDbxnAC2sd15jAFplms6cOc4HH1EfcgKQ86Vs2te0Sx+iuES+ks0sS2PxaiNd4J3VZbcQg4Ofv6
BlmnoPRCQYdIYpE/xBjpIH3daxLrDFsIf8AWVNJehV1fScnuSDGAcxVRdxEwaKXUK1dWNCrL5T56
kpRwiG9oI6zMdsX9cno7oFlf+g30CHREhp7nTti9OoOrZmDENBSle+Knbd/ouEU9lqpe9ZnTuULM
rIY10E4ItlCf5GYck8GeKq35pkaV7RMntKs3Vbyv5oiw+0Y+agycwOnTLBSi0f/G7+FGArU058Fq
cyp/LeEp//ySL/e1o3lfwPojIP/5CUfAajXFvhMXkd+HHf4uSxlVVq5xra3qQ76B/rcUrw+JjbJA
Dit6vgdAKoiKStV04yxjhtqWzhwWd/Yf3bDVbpPS/uOO2Vvuj5s0oigXl2vKW0n+pwoieHiUPeco
dHTX8wGY5UtChFsSNVEiFhgaMD1awRF+nl+2rcan12AZlDm0nGXODPxrwa3rMvDtFyKxiItXcrXW
gkP0lMGcGxlX+pmQArnTuxXBNJnnVKV106FRC35vnQJGvbiGCRymbYDfMTlsKyDhFwNfye1DlOFF
EV62CuDiECtvKhK16N0j4r50x/Xi0C6hDF4PY/gZK6AJPsyH3wNHYpmwATjzGcVL1LEZh815+NyK
Kk1yKQzAeYSBWHe91ItGwl/5cCYXdc1iE16tMwrvUTexl5Sa5U/UCpszgMOHiJ+sIR7YHTrop2pu
wtzb7aOg5lg6pWi/635m+4fdVn1C46qPm/Laymm08eUsQ910I0UYOFLOkvSieSZaIi9e6rkTenIw
GQbjpMcigpS3QP1OuxVn0e+dNaDq/vzedVuvsBNH8B0qYaKwvPNGCsNSFuvk9RI3cq5Rk91uaeRF
oeMkWJouu+Pu8EJv70Y+vwTioYK+iAOjaxlih3l1VJCAo/3dy80mR4/LPhtN/8cYkYBy9TXLBj2D
+wju5dQcjcOU+fJ0iubnJ3mdgmS8Riz2IpYEAS074OUCnBJY4TM20DjP9MISnOPsajfKCTytPodo
2W+AOgIn/ZYXnSucsPe6AHfswJyXP+AnK1bZk4LNrgKXFNfMhEbExE5PYfPj3jG9m1l1W+m9SbT8
99pkW1jl6ysGtJr7rb3MLVBoiX+2wFpjwqR3Kbq/Th9bxLdrx2n6qwWVKCM+wAuMiFbEnYRw9y2U
8OCzV7ii4ltIEwAeUFD55VbGhH4e6g4gKWkHKr8sSp6oA2fFxtivxbTicqslJ/bqzb4VzvuTR2Dl
mSgh106EYlkv2o5iscFBNcrNoBVHp4tUrMNT9JGTO1B/tHtn8tfv+GoDCTY9SZ1NX/NRr/1C+Vqi
eQQIamz8fEL5zsQ7PAW4PLisTsVmiDDMVNiocOPjfcmFmBbnHuQSsbz2T3VVCwRjf4dqIqTSb3oJ
ajOEPFso+66/n5ehdAuAdCXYTEQPV5IJsPNHR406de4sc2udPWi3pP86ieXzn/XiEEUAjTTm4NZz
R3ytlFQN4opramb1/3j9+j/B0j2wZjIc6OJUkRMmIkmvo+ijr3RUI1VXXwA68ZD1Jt2MZbwKvsfQ
mimxmRTjoAvoveikgIzukK661iJwP0WEodMv9PxAK2XBTBEr3Im6vFt4f8LY25Ks9VJD2mEvrWRE
9F1AiyVvkDm0oxEtLAuKdSZnBT/9e6yeOrNDGvJBi1BTu6OPAIDdtW2v7AgcnQMAKwGuM6mV7W0M
9nbgyDYdIAUVxIgzTmeAm5I9O8CmG93a8wyfMZjlcvdqPwFphV3moqqbl2JA/EsRMdgIy5KHoDS0
B6dSr3SZIyzdjedg7Ci1oNS8n6xUIEdBj387esTH6rtmg44t1cmfvpdFH4o5TbUmMnD9MY6y0o80
9V0n7SLOhUgh9EjVf8qmV8s+xwvDz46mpSzfVWqnzeLTe8eB9CqSNAR6/u/t96b5MmbS8OymWd8g
PHnKGwGDzKXjYTs1DPWL0wzqSsu/O5hfgh8JkGs7PjZi0LI6T4yGwa1oCvVIqgFUP+lqJKLFNJex
Js8WXpg3Of5MWcQT0UX+/pGOnSKsel2ZpKsfOyR/pVmaVmh9R9kbTgCqsmXrD0f+MNndkkTVV0uk
LpCcEBGDCElmLXyAcaiNiH2qXWkrQY4Ma6coTBhFouC+VA8F+mKV8jigm5iSDMZOqMGUgh1wEaWi
bBuwciUpxZZ7Oh3hWWtCFOCVhBlBFkpDwU9WDKEL3R9YBuf/6FcKr61Q1LaMnZHl4MynmYfZuJnF
DfNsLnp6xZlNeu3FjFE8TOvvqOkvsX3K9ai71C1Au7DyQB72OhIBwQSgd16GA/TkwYuIKWSvzx3H
kC9w9QPv3WIlTyxeXQ37T12685Ov+O6MO8pquneYrD2DiZ5MYIsMvtCBkzatEs2qhncZWFttQ38b
LB5NPMhoYj0qck8cIxaKGlIpkEJiqP0aLLFYziY3xbeF/erES1+KtTwgiSHJgsxDTS4ojw24Oip9
iv9S9VDAE+LQW3HKyJltSo8SY9dJLuLxxPUxuaicHf8frpK46ZB2odX1LrzwyCFMJiWJhEFIBPpL
SLvmnLd8oFGwz0DDSN/ZflWfeElNS4YCyPoBpVsm3dYLLv6f/MNpW6/hCD+FXNCLvjKoEw75Ix97
ysgUwtGDfh/6PHWsX6j/dMovdX7/Fq6ss0UXLx9DtsZqx4s7i0BBIH6wWXxT6zirM/C25seydksW
6Lni6fn24fT4Ut58hW3NthVbbqAs+NjQ+QP1DMrRRLNYqgHcmgnqbvBcidSxsmrbQUERicxFMv5k
ZdsT8FixODe9YG9CN2LsMlfk4AgMYWsCIvj5nOXzktEGdExIprl08hvkdb6lou0nLnKqF50bKeaW
h7MsiMLgG/PphkS8TaIJh1qNbWb9fYtlqxSENy7ZEt8H65EvcjPAz0VBD+68xk30yaONkTS1drB+
fOlTkFuTxLWHv19JThZ7Gf0xKV3omUy1EJyEScwH/fj5pBW9o2jeMs5iwxtWzxM/oBiv9IuAwL0p
mcTLEpVTeP34TAExSDaznnlUkvFiqp85qwfIgX4r8A6lpwPkbR4L5vpjlZV9/+6hxhV4Tl3mizOF
FdFRbTmKN0XP2F8pqd/uusnNqT/pbsXgEfOyQ7PodX6ip8AYC9zwhBVw04VbTFRJrC2CD5ndK4Mx
NN+ap/SHbxG0VZL8sPTJ/LjRwa6mEJDBOdvFxfICCkH8dQC2Q3lzNVgfFU9Dxs0MfQ4sAZYDC8Tf
9RchwPyZPkpmITmbDzeMVpJbqa8MQUgrfEVTQgxa8BLdYbmkazEPLQkFTGFcX5M6Vu/M8YMA61um
Dlaj9lBre9jIhAZX+7gk3X48z72of+jsY9B1oSzbd4zgFIwU0xcfGv53YgjQTkq/MFbtYO4qLpzl
8TFLhSeQugprHWr3rhyh8gjc6YXXMW6DKCHlmFpPeCOPw2BuPSqO5bQlYYeaFFKZ2MbtAE25qBS1
m1viXtNC965H33jdjx/5eivDhnOMK3A6UrRewTq0plX+o30Dod8NoNWLQ0x1qTf245OFvUOfcfih
wg9Ds0Aty4uVAeGwRKQ7f1RrYWL4Fj5iMRzH1x37sbU3e+mFUdWdmjeGk1zdthzzpbuQQMtXmxvg
ybrtk8Q36VHL9hnjAIp19LftsuZguAOtd19lb7uWEn2XYQ0pOe2nzLkf8zCONzST6HZR5iYvWAEd
LgvHbPFcP7kCnE19/FODyHCLRne+AYWU+64uTNVa7LPk0NqWs+mECq878njP1KTMUOrj+qE43/m9
XdGsdAI88g5v8KkbMVRNW3WMv/O6pi2jhRUtaUFJFgn34hNwy+zlJfF1D1i6POFEGdYpdeuI8RQI
a7v1jYolGO2hFEm/quQA0Ipx/p/K806EiipgTa+NDWoHdKmF5+FW1LVvHZcr8on2lUXSlK428+2U
KpEbDYUzzleJQMTZyF/QUVa5DUdjnrqlt8YxXOi0wBY54N2dGfXWG4MaWteDz9C+DpR+8y8pq9H+
x1iZjS2t2aspTTQQ7ihGwNiGqsmXsVdROuyzO10BO5gVBRScoF1WeXp9jJsZSzCfvOF5wxBUui84
67keFNGRkUPBX+WBKBdCXr0Ze/nHkE486TV5O6OO2KpRD3LLEZfHr3D6ao563uTQvi0kzW+K5NNK
xRph7vi66tPKr/NLv8XKtuQrZyrTAxMhywRiWFcm2tIlyriWN6UKnUO9vWsvbb5k0udcf9EnLU3q
2SXjGotxKSFxvG7nrQXgiPAhTvoj8ot9VSPolO0OP12pEBaIYASz0l4QvwvSHV3i/gNICu5Oy0Ez
3PQAsS3WSVTwtiBVXYcj1s8ZmI8TViejC9ZG2cuAlip2C7QMtngTSj/l/zatLiISvtStGTT1eSXX
lMRYW2jvMtVL1EhFWuW8hkMbxicNr34zWtx433HSgYtFt5EC+JDIpdXJULUYRdja7F8DlGMowoC4
qXM6eTqv2DKou4Nx5e2QpbxIC+SO+HEfNueZPPJq8octxbUr2wvYBv12nhJFlAtlD/yZ4sOVKE/+
2qy7TP14IhDxFIrrPSAgOo2xPELA7iooV4COUnwBjCIVpiK5sV/SJk3yxeTntlkngSCDz9TJsGCX
JEya7Fy6+euYmAh24LTa2PZdVCt4tZMyDUG5T/r0bZi//6wurApG+fg+HYoXMLqnLc+SJm2Ut7Ri
OIVts/k4x2+KcdcPYX44fOtKHNenASqlPmbS2y5RizKS/PbyRy6Rbpd7gNW++e5ZwVssrCasfEuW
WTujSHdrH0XTY1kv+cTWdhyxkgWvAFMmmVzd9TUa2jUkO54PA9XNY9IEhZaMMa9ZcI2i8f2NQlm4
8+DeMzdYjWPLUR/SVl4E3/WwF3HG4RS1118z//wvhO6yawYtLC5aKIZNEwGDa+tp56t8jZbCZ49G
uLKUGpeo3hfhIMhpSOZCQ/EpPuC0TorWDllEng3YeZ7/UvjEX6MUIkDHhZIGZ4DR8xsvdO2291uC
61xktvaNVSdGwpxKBEM+FtvyPte50wNzNc4FNaJSnnWPXVbCb5SX0RLGfiEA1fjjrI3V//JPRuDR
RYZOssMBD2mELwkBV6JQj+9v3L1/gR+drUnxC22JyJqYYjU1lx+zw5DuoKswgaKQHXA5QH4qQfvw
jjW6zg2/ad4AyZ5kfIQRL/8mmuuGSPvD8GwTWeJcQ12GAwfY3b2y0FsWcApnJ1WdOXAUIuabkTBu
GGyZ9O778Vzqel1FE4OBFyZfwKffHwHz+/g1SvRG0fL7CQj5OZXcKAXfYKxEpYixaGxJnXvqDDya
g7XVUpfyA4M9l5KcqHd2bv+kEv8HI4u/NW14AHupFfFysT4CVynY459Iw5IXPBWXnPisK8XguidX
iGSFBJn0kjMKqBjMrlzBdawN30TNF7IoqT2/OFqmSTAGp1hf55i7E8bNnDUOCAyFdMIhMoLRhdpM
mHweNO2ORR6kZ+K++XKmc5bF5B7lzu1t5JCDj68jr+OYMSqoIfb71V5pABBpU99SE1FXUxAzSouw
DFRBlfOISCJtWYrZ4rIzgjYeXE458rJSEqdFv5ZT92Crq6itg3Gk3O2+vlYw4L/tWWqxxdzEGev4
Y+5BIS9StN9dDv1LrEoi32WwTc1vNuDb2XBbtSV3dqpYr8NyXJR43f/9QLaGly3ysXz4rJQRQBaE
ESrj3MhVEPqF1o5cPNYJYCJYq8wgsK+hHBcKYDxtAtj2Z8PqwTJ+5LfhQmT8UapLhwG57lK/dL3b
8YNVtiOQDzkKFDGTKjnztYOJFZokQxcMZ8T7vkq9LOO1DJXHnqWtCsgFHtFMezF4mbkawayw/ch0
I8FJNVrWbyoPA7HX6r7524/YN7PMzOUuTFL5L4ooWBY/Fulflyep2cciGXCIITCMgX3r45TY51Ak
nLPS0EqomTiPDfd1Vkd1XDAB2lopNQQuBXsGR578JoETn4dEypKi702IZJyAfnaFiK9R6e202KmI
UFBXdyId1XldHDcswak+bP8pPY+6PWW14gB5OTxDYJ+OiWrW8evWdX0DdyVYDVnSr23eUjd5mCBd
KioeW0lAfVBkfFnJfSGb4U/Dd4Qws9dD37SYrmPfU83NniQW/3h5Pst0ak5b7/TgA4h3w6Tuf/R7
0jY6nRJ6/Q8uHbeSyGY9ME0xLfajB1vSK7cv3PVgx0i8tyBFro27zXhMfEV+gWDsC/U/us14RuKm
37S8+Tbwcd8BdjDtqAUIKL9SaJ7w1cEzlHX6G0tkrF+5fukJtUpL/mg/uvlQufmN4g8te1iwvmWa
pyVELUusdZ++J/jeaSu2QXEh4RSdyOBXYZ/6Xz7GLFg4ozybZTPOaz1yP/Lbvhid7JeLAxBEJJQ9
GJnyV1bEkXn5GIumVh3Ct0vDMuAmHmibxGy7u9w+sQbNjDte8kNVpeVhTwosKXZAmCMVnCxouXkU
Sx/UNbhwWSgFcGEOke6yhKpTFD7shjeJLB3QEIIxSEH9dcoO/E39XpzkoCwq/IffK2yxhxG760XR
s3b+T70lp3VBWhbjhL0oB1H/zH598pZmuX9XcdEGW4lOD/eERLH5LJXWmUXixCPIZiwCDYfawxQ5
3A6zccmrgxtEgbqV1ZU+HLFvcqLpgc6Isq8mIxsib0eIEPPpWq5aaTjzudG5sQVwSL/KMrkuojNr
04K9FERTUfOEAZFDwJbwwdcsY3NgjQ2QWj5BDQ4GYv0H4txKz0AcXznKJuMFHHx4GCdWaKjsBgpH
yYSI3zYppC02ojO9WrA8wAg3Eh6Nl9RuwQQmd7Fi7mCAA1n24zdAkK0JQwRrg6Qvhvql1F+Q42Y3
QzG1biRnFFKM09RZMj6d11RvKUX9cI4xR9ZL1w1zB2yBhNH0oStBUiBSlpOk82SJ/cJkvX4cTUSE
ijFrJPPf8fDVWgbPwcE/FNgMT/G7Hltbp1U95QmdB3o5D/1Zsrn2/XaA8asJa0Df0dPOWiZsq6I5
4FHQ+C2eEV/UxjnVHYN1puN0vJR3EhBL7h9TkQGama7dDOuy59WLQyRVO8h4+dHLX28gc8qqDITF
bwfAHHtqJ/LidB1BvbIL6Ur15caN/rnjOcQ43MuFT4RuY+PmoPlrKRrJNX0XEKDY0FEvIuAZfjve
ZKr0H5OpxqsMD5sJPjPoMYuINwrh5ERAHaXGA7kZNqRPuXE2K/Rz/wQWj50oR/L2xx7DTMUFFKTx
uKRjppf6W/eZ9F05vz9chkbjNKf9ZkBzmCipBNVl6xcyula0GEhnVLHfCLW5PfY99JfrfO6Lakrx
TbUItmMLcXTX1OjpnrJDAuW90ISUoPmM6HHcDmmHAjmT3db9rjgGbETbMp3Vnn7qVhAwKzP6Azfr
g9ZFtbIyKLbi1IaraGg1Ol76BtAjqi1L/hjJMrK8QplHD75WVVW75hu1eBGV5rA+LvzBeJh1Zhk8
hafTbiinibV/ox8lWBjJb5a/tATotbHEfGAXK6kXXzffArDlqpTYuwimb4oLL9eQHEZcejRAq836
GfWUOOb1SkE7mlMXo7xiyX3oJFvoD540rXzbfVUAR/bWZNiNXvVlL3AfH7SqqNIWNEEkGfQ8gKwu
iaU9GzQIqCfCWHyp/o/4Ze4tJ5nz/kxRIwK8gWiypAezU+mJ2uSnZck2hkTgyKWVTNgwmpHSbwBh
O7HblWNcInM6iBdeIaZdWkA1GgBhRZfTUH1NUMbIX+WdNkGkIGXgd/18lz1KIoLUi+nXJG3qWCkM
0YstXYPZEGhRwWn6cclsMJJhlMCeA1DxoxpUJY327+ZrMZ/O8dJMpU+93ifPgDAkdgh+V+ZsLpY+
EJAA6GtQEwFzDv3mFa1n1R+QSd/9LIG1lqoOs98ALWI9fClbGEwT0Rk91w2q8bhk/+GLGbSkeYFT
j4HqfcwN7uPYljp5nsLtuoWmXgq5Z/dccLbbOfryET0L7BGGWMRyzJUiNLTmvR8qstHWpOKHmXDp
uh9SkOTebxPV898b0HCvUc+cU1iGHR+dqn596HickpEOdcoem5JfEyL5GNaU8qMEDsSrcjrZR89E
ITEj26eNsVMuj7i3rlHxg3rlriM5xF2OPbJgtQp+v2IsWEN6zw6o9ZptPNsotzfBSx9hu24drpma
b8MXJVeeI+kRwckEtZBPnZDKF3IQAS3KrXPvRWjRYoaov4yWZSOc9rWjotfDTtA975V+gcJjxGOE
8SrS0ClZiO+iSgFCeh0kN+dhNQZwndWFJsBTqXUqQJEHTmN2Qet79vrmAfR5hU0Fb2XcAwxT5xfy
EvAAxT7SlKJBssIEhzlDUdyTkxXnL0ElLfegaewgTPvfN5+XQ1CxJpC0+wnMU4JbsyNjrSq6BuGx
eotaHl7xVfJ16T4LHCVog32XnG4CDimp76eMIT6Q1PcyVWQoaMPtgv7VL8qeE+FF4p1ZkIm27i0D
mA+3w9on3co7ONqaXBpQoeIx1TxFtmzHsTpQWOsax0VDPtnoS2EwDxnbaFEnd9iXsIe9o3mFFpCC
MAZwb5bmGrikzekAiIL1BMxkVLjLwhU/zn/4Cer4cCKavjT9CtWQFHCDM2if839EzSJSuX4i2jEW
UMiXTXVCqbMVvDdycCFja9nej8IzKzbUQvsKDnVTKYmr+3ODbzzPnbu8jZp+dQOA8tA7+uqTt/Q0
q+DsNhJc8uwuSTnpi65Sk0UA+V+R7+ocrjSHIp00JbLbPRjwYwtfxrv6uzEoQoTy4LRtbO3p4Pa6
haN0m1PpVe7581smU3SRP8357XIjLsJwChrm2gou+RlpPOzl69O9qgSuU0MUHIm5GNV8ZKiDFIVX
6KvVpoy4OOTt5FloR1WZ/Df7JIEhnqgOil2Y22l+OipIvwm2a6pPFYMw0m2iCoXMbo0lCvuN/Jj1
Qp0gzmzzuLBY2t5nRL9xuqDwL4F7Hrvo6aynkOY5e3uosbFieYDfKLoJoyRB6ur+2pbQbGNiqDsb
GwS2UfGQXwSQdh8MGJZkLq3oWB3apx1Jrzn3nhZtxpVlwS2biKM3dr1iGbiaTb15jE+9atHG9Vax
USJRcYbH9x6kCb37DWhVBgBCoUjkL746bpF5YHQBYOzJW8BMKu2XtHFZbjX9NlHegfIUKBgBjIrx
4Lss5Ve8ZmA8eaeH4dgKe91C6sRceQXZrNzRHvaszmFeAb5zkHKVI3mbgmeaNQTQFac2vQFsgqz3
Dq8YOYViHAVO7VRo3g3o2Yq41+F2iJUbIE6Gqzl/g4bY31M7zD7Blr1zm30s8hAbpDAtIX8ObkEw
sV8EfX7GBlyxMzAZbmDFhx9HeVOSw0UpzmOw6KmFT9DqjqpsyE4fnmjv9E3GXnuMZLnkV2X7OU1T
VoSHGpuaun6isfe4//IZflWVwBJbvNbSBSSGMkv/raKyZ+GvqpHogq4pzbayorEqo5G03ghLvLMS
2sHuY9ghLuJUmWaiBbHRmoYoRPV4nVhLwESl0BRLQo+BxzhrkuPoTC8yrW8099x97HB4QF/1/kR1
det0BU5EqifYkDLvu7WHIzgAwDCiZsHkY6L3QJ7kGmM4YwuPaW/P96HJkd/bOx7bEPZVMtHGP1Px
3+kP5H6SVOeyDoULeGMApyWIFohU7YDYBdEmiDvHEzDB6osfa46stqqADEDv/7l7Jty9SW2kxPyy
EsMzZeoMDhqP2/hhpFENYolnj0jYbsSJUGPKuoBpg7OmEJ1Ve8woqyLcmKZcoePZ4vfpKhhaawh5
XUbny5ILflcD3puwQo15rwRwx4c6Mm0JEzMRjMZ2gRqYZhp0b/rF256Z6aT/VYqDRJtRIi9tcndi
CgdL9gknFcC5QNmIC/6jU7cHBxP4RR/npKfHt4QiKqjSlA3Cr8fnsat0687d5aGZ2mk/sLb6ehdu
fVp8o3OxEYZhH/Cu/CJBopDMHwKTYLH6D6vEP6MNNUV2MFlPbGDnGSrXsBzH7JqMEv+Yw6v59k6A
RtU3/+oP9roq/gW1YlffO0SfL+u0DEq255QChNwNCOWrxGjK7GbpQ2UQN/8PU8/gy/C9p2wE4/a1
qJeozzgRFcGeX2/vWqFoegw4xONPqarDVSsaOxZOHsuQqUWWgs80JjLMa4gwVrgMyjVdKtgEgU8x
mwC7HK5KCjNy0GPamdHfVAjiA3HWHOgtg4otcdDbgGp7C73nI2qyWljcCuzzshlSmUYp/2a8svkf
b5ulTMRRUUoUho2g/Uqw8s24ZVDtX0NUpTOIPhmzVn39LgibUMs0Q3NI3JvXXJjE+DLSuJB7cs7A
6kJsKqDfzjX5ZRmAmXM1jCRkRgHOSWIsApPhs8mZMDnhAflAKgm+LY57eyYH+sl2YWmf96VLyYYc
murKvJ/rTN1F+m8/deaqK6ucHnpX+ouxUq7U2UaCMGVYAaWDFdC8qB8cb+vZSpA9JkBLViaibC5F
weoUAn034WVt28P9wBer8FECuzzWOJQ++nDghny4pHxQ/hYybdDMH1CK98htzZfUY32lwhAk6kbu
gPur9OzU6bWOW7hvK+Fwy19Z9bzTIP5erHudlBqDgzV2tw8Z9da1xgPe0X0HkUn3V8XibsQOU1V5
QwX7IqcBEYFTGP9Vp09KYpYfBaQceoJgeKQXHO+XUodtKCTKCEb1+wWQUD1U6jwy+V5cay86s/xo
6Y/QMQ3db3GHqwvk29HOobwPjcYsM//HMF8ek95dfPXxSZRvLAD3/KmtKXJRPVzRx+/GQWvEJrJ3
zGvWAzVRJsglxSM89IyhFulZbnR51uoZHeu2AiEj82FrCbpYleGM+3B4ICQiMYqmgUAIoAl2DrnC
rkkjBKPp6sNxKdvfiA7gpg/LzvyfRbpuy3EpcNNqH2ImZQRUnhKZSbVBRlkOObmhG6a5YoBUASPu
IqYtPUHYqLRu4+ma2RD1ZdEAR4swBWZDEca51599Yj+9n7n880ekFcbIaYKc3S4s31BB6Yu+h8bZ
2ldS3ZAJXzac1dS3J+u8ObLiSzfaELxF77s4YBWkkpxw7YbKPr4RD4AbhjDhDfULwxaH44cgyTb/
yau6wlX6pII8jKq1dG1X+Xpz7qxqhLKqWS1p1GHVuyMcJXtqpyKwAAoS8Poit3BcOYBu5AN8TEzR
PX524NtXYgDP6p4cHZ85Xd2ZGIAm8+5heuHZFgqbKEo6922VPd5a9Op0nctNb9aBa+nWUVB26Kzr
185dFw0ukUUYgtR7FuP/w99Dtu9GD39EuP5Gz2jiTBeXRzfsl1HJSeDuN9YO3kDmQJFoAApPe/Pc
y+AMQLBK/67Pi9wJoGFudpmzoyKbz7xUWR38T+Jt6yFJ8/+syu7sLYK+0AkjvMOMNKyFnfZpx/es
2zm9DBtgj3xLXzUDQrsBeNIoyBN4Z8udjHh/N0Eej5NjyxdQ3tmRdb41xp629MKRtLpCvL+l+pXG
M9rZL+XFgr5wkG/qm9pDTFzpXnXQBN9t5IyT0cOvUggzQdS9tIdEgOnPQvI5RdS3/gM7TnEHmigV
4ESi61VCnaXtwXPSCbePu+BVOg4WHwtCyAxxO5srPHNMaBGz/EUR+HM5I/xTy0IzmN0VzQoCr3L8
8QEE3GXXMwCFOGkoD+PzXVVCaynb0oxKDrzoD4rA572ujLl55SQP5+z3qeotr/DEqvC2uaczuect
TZ9HfsU3+LlUkJk4qn8J2pHCFw9WUTkzgdwQqCDSIQqBP3I887kdACcuu2CF0a4IPgLwPnossuJD
L0+7yAgUZ/nrCeib/DL6AUulkIE3XNVSrHCweWcqnynLCSTRG9KNslS8GNQVNz+qYC369mx459Kl
48gllizKoN7az78QiG/JpPJoMSZ3cgTOEgjC7rtydGjesht43y1uca8XOf5+HhI94DkEyFYKZsRn
ABXlaZ0LI5IiOmt7ekUC19Ra7cvJSRLcHgse3RnwGcQRv+M81cnyYkhHRDVXwkah2ibqDBAI5N60
FSeTA1bLqj/ZE8eXtLX1EEctJFTMIMv0rx7xKPlMfSXd3p2jJT0JIaKM40WIooTpZAIZ1TjVG4Ka
vO0vbS14eA+6tpSD8od5rDosSVbMNZao0fPUndF+zfmXqL5qd5MrEOHFQ8Ly8ovoCv2WBjX9VexW
0a5Ws6QjwWL3ZTUya9dOfUEDckxugApVb1+TRTeg+SC6/xJTiZXMBrmCbRbZcl3oM2lWIqgU0rrE
gHBQP/qMwaoMmKgDsT74Xs39d/3JOw5ESQFSQDo6H/sSmGlpoxKvSJFruqVanC65T08B3msDn2eh
OB1nUyM3IRApdifd9JUrHprSh1FEuUe2xOPy23FxTXX7qM/SK+jQSvRMYpaCdL0XDB9lhAf4aYzI
U+QVYjGJ1fD0JQMnCid59rHIncP4kovKJvnQqJ0cGCaRJOqsuSclpbzA2D7HzIiK4Hekbnscz2t4
RJAxVCpALuVc97YkHakYp32SzjoPdzTUZ6hWkF2hK3qvFUUCy2ExnuKNGS+/hSTFicsywUO2/WtM
GEGjD8QPXsGa2/UICW0GCXEzfw1bq0LWVUuSWVmdLa+s6KKnK+f998xKW0Nb0zbKIKyTEKHRkX7v
YiPGmy0Cyy9g0tFPJ10Ukq/KNroEv6PByO+Z2k+VG+Xbmt6Ds1XdqEBmeqg/wbdUzJ17km9dDq2X
z8eRqKBHzUEejwMqPgZ1mfdEp/4x4ngh3Iz1Q1e1Suc50YrRxYwFMlqASgv1poqzFeckR1DwGawP
k3I6SkJsxLd1ViTMXspZMCyT0lWW+32GFRASHtq92OLNxJE0grHxrknzp69rT8ka8kP5cski5t1+
jQ5eRHJntZ+4UxfsDB0hOyyi3l0MGgtaxVblJcfyT5QVrh3RZiUPLrJhF3iqMF7y1hXOhoU1Sk5n
k+IjIySzOieQRRa1g4Wm36D5srrvqkmBVTmtGyj0Lnk9v4eAmeF6nmyGxEGTRCF7icct3WSaTopL
QvNFKRd6iZ7OK7mKr8ayT9rZWtZVVkwFJbbbenfFQnUSugFTrHanNSV0l7/BxAMVc6AGnYS7U2+d
e/G5RhqIeDVY+tQanGbVP0NzDt5hypPJ3FAsxtdrEnK3Bh5uWmDieY1j7nT2ZqZUI3H8BcAR8y/N
GmlYJfT1pQ28S8oqzfE4SQ0V8Gj4ie0g/m7Ra23lEXBOLRVCMg1sMLyx9zgLxn6ddRkgiiZ/AAHq
6TLYrDWGZAeVvss3fG0Gn5OfxY4y5GrhHXOxjzfY+rTRMDBTouAbgVomOklQuvMkwLjsp6gomwXp
bHqqTkShMEed0qXwYXIRdjbg55okLGpzIOadc0B417BIHVQYVjWzIh7HZM0E17PAYr+lhSEzsJB2
XQJJ86/3wT/vPEl+90Vook7mLuKssd2UAqqvQCLHU5MFkdCKLcMZ0sj9hk73nwoZq4pqAt21ZX7O
HNZUceZLiguJFIaQV45WJtO9yMrIhvWBE3mpybE1Z3B3R9OpViOPjwoy90u6Gs23VxwcEFRFqXBn
Ztc3sdGz257BqzlePAfabZUl2INTlXqVUTVpm531UsBJ8cs9gdayqHgJ382MDl3hG9Au/rpQRSlz
A8DsTrg5TtF6rBLmY6oBuPBQhdx78udSwX5LWsO5y0ZEdVgZubRkF0/5/u8DdL51MNaBtjP/s1wm
aget7SJPUaa7fNwLWjzsfQh1WdLdOfONQt2qJwbx2XQBQONt7UfVdlQl1fm1CLswvyc/YKoW/X8X
xNaJt6jSl60crpoqjbOoZIgh/krwEe0P2nHGLqGLlBtUiRHDIvpaJbdmwJRTNFg8wmxhsIqUFHdZ
sn/AG7pvHmRNHGupzc3ZMygkJY0ACLdFbJ/1F1u9o1o9y2FhkEHqX3sTjKJvytiRGR20UiluiDHo
FE7YTM+H/G0bxalZGlCBeRzLHX1a2+bv+Fh2Sb34dxUicB7k+9/j9FCS84uK+lpkoh8Zcn5PeFb/
LzyOYPv1f/Yhq57hgVzyXHjXGRXdmq1owttPMuVgj6zSypkKYCljPfnA7s5d7/jrEG5BeQyZWvHy
MjPCSS8pLEJhXPbN7CE/zOftpIqo4ARGKaIYV3zMG6jRDGCE1vaEgwlNqjOZ3nt9zOvyhrLtrSnR
tHPF8N3JbLvdIMj1Ocg8KoQaHgX7MFFtpBThUa0nxLKDrmO81xqGb+gBw5lUwLozo/KvguGDE9vM
axIFmTepF9coqWCzEm8VHXedpnCbW+MYLJNq0kSjhvxr7zV1HV+bFhuvOmwfaYbQVWTr/kWGEVIh
6L2hAKBFzPBu+tHocoJD47kKEicX7VXN7DOdNY67tnolrnPWI8MMCtFUWu6Bd145elTud15Csn9x
s5O7jUfa97oPv56+wKmec8EOcMN3JdUESccSuNnLSPB3HRqjKvp5KUw2BrALi0bCA+6mzgGeH3oI
hjnfOUMTvtMK//L7geIYAT4orq5uZ3cYdSTeOVglEJEFDDDTnNnrAQJ7T5yBtU0KXrYM6kMm75Tj
GoXIC5zsnp1uYcRwpSXGO+SCynMkgDzuiWVtJ7H9vDY8eh0O24gfk4rwyiEAPNLmjodhFH7MTfnn
KVrnFVSID2hlo/i9MiqbtDI875B1NhAgVms1cDtsqOeSgYsHqgWd7RcfBK6o80J6w+QeaZYivwDT
hLfhgVe7wqHVhQlX0JNgDH16o21cxUnq5WNccYXJhnGC3SQ937U9rAbm26HwGbAm30Eg/8xe8c9C
A0pYwSnxQYU6sEbZUqSPpaHdM0/U003D6bs/EYWcElAbnx1PGOFWHhin46KIAPWnmVxlmyaOuIkW
YDCw49h3mEw3tatFbCGETkz4bp3YwfhtCHcHUP+FypiUbFlcDLrRWyvPu2skTIhHlSiYrGyuXrmx
AM2A5nXPzzcFqH696SO+ENaoua81JAOIjPOPuRuIQ95LTMv1ftM+o18aXbywZTKleov+/mc1H6Gd
cOjfAKs4vHhc8muc6vWhKFPzrqC/eO6W/Yc9TQSWiETBNVjEbs5Owrq0wNPXZ2JRzG5aMD2Xwlcr
fc/yUZGEPNXyRFGwkYCmjxLun2vnpUEPlp1nl8e0xEiO1gvhBbJ47GQSahV1BHWhgbV4WFirUQdh
aWrXa1E1u4rRaeGXxFqKKDVuM/sxvTDrH56csP5uZUtVDFVZD5GZMIfBBP8B+QftLGLK/Vx/XItm
rqvgYGGoWAxRu5yWD+Rg2K9Ul7r2W0mGch9TsZjbo4Rn/0DEhyvhArvxOIOHhyfLJNb7HK9JJuDn
MztjpsrFqk/cqTj9sXbvIlQx6BzExnK+a5iQE79fgOMeHiBQi1u+9XKgsRlsfG+eatZkTCACIKL1
3KOrUmd0TOv4bcrTbbGM9z5VysDg6BoV/JEQy1V4rNgpfu7Z97/+XpeaLHIjGNj9vXnMFU0BG0R5
AEj6K0Nj29elEOd/gWPda07ioJRr8BOZkc5UxojGb3JOJAh8XB+mjxxmxibw2vaCcGFdrUJZxngK
AhgSBUFPFyEjTL8eQDbWJdHGiqi1mKZ7I8Q1vz2nl33QnBj+gCY7MhKtsqSa1BYtASPw/ufYR9jC
3OVnEJy7RAABEuWZqmTu/N9/uJltwEDDvEJtt+IWmP9g8xISji6j9dTaWeQIfujRL/YTbTSUCm1G
yxAl80PU2ISbb7j430TTmBeOizU2LnepWETujSJt66Z6H8ghCjXHRetlFheP/2RRu7XNXeeDp0vZ
EqAmbgYMAqlilmuR3xDtmQaUvtcopJjp3G5Z/XMPLs6VX0PiT6WOYRsL8u3foXfMGC11bw0bSm35
fLJcCE+bWLREw3alxka353o66WgVO8yIabM6NJYAHMK1Via9Hf01Uv3IvJZbUS7daKhAFRi0kKZC
4hZfZ1cxLKjR7mpd+vQ7V3EV8AAx+fGASVN9j+kE8+bTxpzpBILIs4qQSs30ca1lK6qaEQ3x8KKJ
vFlctExkK0NG2HWAcJ7kzQgvl76Z9YKX6Nj+6rmPTkqpNwEupFtym5t17pFb73VDF7+5N4JRg6zi
UQjWdmSIb7imuPsix9obut4IKRT8OZnuUTOEXHbqdP54RBgbPN9sAm2heDX4cmk/IK9ooYHbEGuD
xfgYuIuQRcRMO1/rzKFZx1yTCNukqAvv0SKi1//yDqJzOW9nCTRcEg7Z9hQrGxDp5UeACB62CTpe
OEmloRiFMGN41zRmOWHExq3lXkre2sGorOZWivpH5TtDjx98iARUjSnVIfzzq96OEfGDNxiELLiV
cYRkIi8qIcy3ohGTNBbLdoqNLxkmHxNokUuyEdRmu3eDg42eKpiOAhuTglEXz7FTM9UkmYSsb4Es
e2ilzohUzgR36czgxs9qNGm7iw0s1eYe34XM3P8eh+bi7Yk23JTCwPXPTjZyT7lWQ68FKArYcga9
tWMC75qz+X6KBE6YM92g8a49yls5torRwNDLbZ8DzeQ+vbgSt6qVgTyZ7bGC2BCDAgLI7JmYoWDh
sMBwRV7YBkoXcI72OQcr0vKIN9/khhhsPiEgZuhLs06wyeHDntm8thPaKB2XcrGUvwcBD66QIjTm
1gPcWRqUVPluoQEFF76WpytA8aPbwAnV6uXbFV3PZ9GbzjSgw3eOe21o8P9W/Kgxsz5jZM8kaDRi
ZxprOOCYzM0b79Lz4varDu0Wl8+CSILhJULnkZo0Wxjboxf2NafXbkFGkksugBJBVcdd0YIYjrWi
f/60ofpC4PwFd6nXTa5clfJA9xlEqJS9VFif6CK+xS8SE7ZEInHp3MKMVq7h3TCRx+N1NYwamFgK
bz6EFEQZkV77CxCV1RgzDTdc9DiPQUFR3EbQkkMm1Ns6VF+IRd5KcyosFaQN1bDaEner4oVpCOsw
bdB2gx3R/a0QswNkyD4FcmYFYDgS+B5mtQ92Af2VISkn/fD93CrR3SjEqWxzEvOIdsL/2FRJUzJW
m6E6RVouptFX1YRkEWG65/BVs/gf90Qs1Hl2Qhwnio0ol18HMpAE4hIRBiuAS535tQpB6ZNBcB7/
+25dkjUVeta4bjSlsnphUn410i9/cAYfGLu5/NIt9R9/3PngXtBX34d00vGNaJGXCj0cmjsQivUz
c64RuN42noTZS9a7LyZJn40xbzWhGk7wRkHhpe8zUBjoMzzvD6/JwJPEH7H/qPrxRRg2ucscfZgq
FZJus9Fm7p5cHdFm2jDiGUH7jzUXBhV+sjQpaFoPtJcnpaw0ehqt1qaicRzByebgEbnJEhZ02+8T
KJesiF88AsDxy3J2h1OD/piJ19W4kUZepe3Od1zo7TRCtwOy/n5qnF12+O3ScK3ZxiR0ErdI1E4y
8W808jr1yQgEegSv5q+3zvyMOI3UZCkGmdvPRrucM+qlm1Sb7w0aZy+7FyHurAEJahGg7vlW2BRb
AHjo5xa+/OM5AaTtU37OiPgkPNRQ6VbXv+wlYosO6KBV4Q5WuFrPXHgFOVSqdEdF1ryIFL3O+xIW
orPuCDivCNqjjWQLnCT25CebzWLkZaoJNCKW13Wgkik3WDT4yGqj1w8bS+XhDFTg14EkUAjaGk99
FsVCo3x9U1xOALUoq+PtOtJZnBNgfvCdECypJuWEnHKvSdnz89+q0QGsgFgFyQcd5UqfvqsOlFPX
1KNW0V/evvjwG6rdWfkVrOqu0i7Tb8qBZ8g5cc2QHzTR2KTWc4CmoudbolvnIDtuRVQp4rw7uCEF
CmxrCklZpL0ciJKu48v+cpfpTDFWIQput495C06ptgp2Z/fiKTEH5Gh+NP6tFwpL2ybZt2yirTPh
SoGrsCDbM8IcqTZZpnJYutqaivCoVkvxb0IgVEUKU/cZzNjOacv2w7t0L0Cu4SDrxPJv2W5v9EAF
+OGvTsIBERIlnog3ngTwMhy5xEL6Q7EjrUi5L+1aYnEro7HKcikvOGGkW6bE75ZmBRf0hSnvuYRB
xxEtjhTusIVgCGWpyEeGeMi3lRXclz9waUqA+G+33YEi/5REBizl9by0B0pYhq5bCfIUFuXZrNBb
C8Ja5/WRLGyodzKk8ti3xS/PBH870727mrcxKsID2HqNIGJ7SNvNkKn003C7nymQicsIDWStc99u
czKlbsb7Z7Wm5I15REkbMgHZX6BefBjPklpiMos0P8tgBdRkgfiVvAQy5hfFOqArDVai4sclqZWM
u2W1Qs1kleqEe6FXqW0I5n2/77gPVkxSOb+wvoMEIkr45osNjS4Hva9n4TrjupH2RZhqz5mA+SvA
k2AsKLK45ZKA2LI3glbB2zt6tjAWYLklzYzEvRNlU3XSLWyJPxk3x818my+iO2nP7el0ai+1MJu+
ZXX7JP+jNM/9M9DmyfjhW+y75SHBMeeIUDsGlURuF03diIC7kkOCyCga8McK50V0VSY/IsOTkoX1
dU+69Ifk2nAEu784lGkHy9opOuNkHlQjX4Kt+lJUbNJ0vfK0vU4VnCCCamQZdoyK6gBhgPxCC1zY
uzDynVKS3Z3jcJmfrus+Gj/MAS2Aals0Fk6q48oRWAg08ihKvAPnXy8B0RW9n/u/86BPfKZPNPD0
48VjRH1XFUXJEH/t+EXVxm6FtvhsREGkdMAv03WG/JyyU8Ts9bdsPb1ofvWamE4HiW8Efo5X6dfn
XZnGvO+Q07NARmIWy6juNvBK6q7Zqc6lKteesTSwsvXZEhr5MgtXqqXjbBhf7EqOfYqr4xQMdZuY
Csc45vVkNwSUqLlIPZUxk3xKu6sP4ynvgJ6KUDFjmFljcl7hn04b4lxkk+ewEsvxqqvdZ/x3/tmo
42/ZeNy0bBkT4fddrC12sBzKr7xYa+0aNNC1MAw6pYkzTkjTAJwdN1vjHE3cVFtuA8Tx6XVSHSL4
FMez234HMUr/vuxGRxSZfASmKx945ZJ9cKAmLikR8YkabDgmUoRrQgZdrBRaETqATwmyYla89aQ/
d/uF86bPno9kU+j/1y+WdM2qStXxTpkV+5qFN5cpT1P1OBkyi/cSF31jd5dOXDvk+6ghmnDE54v6
RsiD8GH72XWZbelyPJbF7TiQeVGgChUYqS0jcaPSqhI3sgCamk8NX3EqTfizI162u0nrYe4TBEc0
R7eS52OSLSySdC+/aQIW2Wyk7h4gFIyAnrZyH4qsTieGZ9M79N+HumrrD0Pfs0F2A1oHMWCXwNVl
N+4LzsfqqHAKvothQaXeGtLYWndMizbj0wxeEQlhmAl7ngODCOLtEBCDYI2TtmEkxjr36FNZiLxO
wIJ2Z7MFwi4fKWJtebAcTiTRoOiwmUyIfBQmQZe2NIwJjLPLDlcsTebtKpIb0VMhjIXbq4ziTcI8
nO+FR9yaTyatz3o7i65nljc2tzcLkKlFU40/vXMufZJEhG3/Fbnc0p/tKTroNhjFzS2k5cXUaFC0
ED0ICw+oGgAfqr8Ct3HByzuVDZ1aBxFVZFmsqgvMor7K9AazXMBSRQk7PceQWYw5ElXpu00NmJ+C
2yiJ+FO8xZuXAchyRtjSRdjMxgHyjYBYyk6IibFLD6odx9wAlq/C/P+uHYRoWOdm/5YzQYpqHQ5M
YzB6nZddPijO5CGWWHc4ifLTSdms/o0iBZAx8np5jP5E5NtNWpDiWbDYR1wfTESNQqLusBy1yWa8
Zz8+a6SPGDpkWKfkOFFP4xLI4HpSaIYDM0FHZzWKpr4T67iBDDcwv57tCDRmUU9akxvHK5HvAalS
wUi3vXx9waJZNChSZfbcK1E2iO5rMPypRBGykzL7mi9xxaTvaQGixmY+BQbjxNI7j4nIurvPDFNw
zs89+sZRGq0n/Lzuqch+H4wk2P0Oy6rZbRq8KFHkFTNjwpOZdyfiLTJKA9K2cAAbVXrgYwz3yUm8
aXYY2ATyFPJqIXLJ+yv5vf6we7GTcqsg0nkRqR52o5dLJ4J0W3XvnpHIlOW6k+fjzSSsl2n/DjP5
Wtqpi/4u24/Oyr6nTF8G66eI7dnbRWKoOHH3i4/o4biQy8LfI8CEHnIY7I2xyYewz7JWCYyWI8tw
2ZJBtcKNi74DwOwTVOMpavYRafbS2NsrTJHpZxGamuHQKGNmVq0LxFj2nRTZtClT636mUyZMM997
KQUPQoviNe1X4spo5tJXnjKzzxkrROnI4sET59oZCK6l8VScvEM/NATnWP1ad01P8ChOvB4PtPov
WJJXW455b6JvhGI920kraOigy9yTbi8zyQs4CwBzCrmdWU+pfAJH8Cu6LTj91XA5b6Vil0WiENwE
TOIEfco49hA0SffxY/lSZ6XlJtmUDIqqxquceEWOCVNDflUDo+YuA3TPQ6b/mtYvA/cBivifz3QP
IGjShdkVHOlfxLmRx47EPCoB6t+/LNLb3FRR+a8+aQ44uFjt6bqEEP125RE4qQIqPIqMVoJRfvK7
7pm9nEg0+OewSnxzbujN86AVemo8BhhMF2ancv38p7u4p6y98+FmZLvp57q7I2ioTnE//YJO2lev
3ZjyJzbJxanSC4NdOWIzToPz1xozOX565jIBr6vRiqgwvb/pGBU5Sy9dHjb+BWzBPgyVroB2SEAW
+4fwlkMDuZa+jivI7ePXCUazMKezlxmqeavW19X387+gpVo+UPbYx+AzfJiobfCW9htxJ3boREN2
Izjm45pCaRY6xcdE+u1y4+UiygCv+pKmchUcQwtaIZn7epNqvYbe4NeHqoCbC0vSl/V0wYkXjJZ6
A40UUBcBQh3V0oD2RdYc5Z/ja1lf7v/5bxTPmwCJCcceG8HA+slapM4+X8esrCqSB8OPQhOzzm8L
xUmftXYoYXhvAr1wtCmB4V861oqlGLEm1YgZxwe2j9fsyU4oAZU+L4SkYm4v5BGFkfNQLzndCexz
rp54D/RxJh4xAj0p9W+MTL491pUjZNqu+XiJcOlZnRgViX40YjvK1SFCybrCMK4Xc3IFZBMpljzO
Znu0joSSYS8+zc2+FOUXWE1Xq4znLmTU7n1IMx9rrW/QXg0M5IyWH94x8vIom7GHqFnvyT/5Rjse
LUuX4MfDQiHW9NFEAzFRhSRJVfTq0sQHSZRhN36H5lyYYbo3tZO/eBPMCoFkRrH/3gu8mxylV9vK
MNtmBVen7cyFqYsi1XuEPu3bGdTY4NW6oWSS5Hk12ZRfy3gfIGs/tOxB7jc3xxkejXMZvTRJi2SX
S8L8L5G9CstaLFFjgkAY1Mo1hAvbmScF0NWNciogy5TAlhrsaSOMsB3SXHrL7BO1/d5koFcqb0QY
yLKe+JQFJ9/8p1+T1z6HFjGbYbzxxhd+V+kgqH5xJ/U1E06neHFoQSj0KweLqIHJ2+eJTXrIPu7/
mY2lUkwJB5Icy1vThEPkE5ALxtMwfsA14VTseoWCuatqXuZPBvSqT/Ef/sO3m5zxnA0Q69pmzNxB
12PFg8qw3mxZJJmaSqrAbsmBwNQ5gMKcDk0tku5rU9SgModAVh9eHynzFd5399/52fgrKwWVtZFm
a7wxCUl4yoKUOL6M5i/VEFW/XJbiGCzFkCtX+oECu5UaPl4OUJsMT6gw1JB73gIDBOtu+daEx65q
Ov/5MrBoU1L34B1yx94Fzvy0DanMLvzaqcTd0nLSLKRVCweU9LmFeCpRS8LsSgEoLMeD1k3lLHev
wq+HwXcceZtu8OpGaATPE0p3Br7oU2ueTj3u9tPVF3/8hMT2M2t2FlIY4Z0gMttatIVA1Z7YjExy
EZUO4uoooXD8Gg99JmmUPJWs+Rr8/iXLZYhOzdAMdDQ5GSBfYA6Mrp2u9mXFdykSwGrkcfiOOKRa
YXzw8ZFPQjbZ9zTt47bJbE8WpCtK4xQETMJDz4J59CCoxxZB3DmpH/QVao2hW8H1jIgz0hCxmgcH
8BxQDRGdjhPVPmuAY640uynMVq4aL79bi9OG6PNEo0N/Fl+Kfq2aeM0TJwcNqFls/SwXzC/lIKf2
opV41X2BxAQZ1/TOqJEggjJolhyZ9/mmeY/0/Q3s5dAqBc3XY3XvoF5JE7riZkVVM+jbrmBcudlT
KbkmGDGkiiEACy7d1gikKD9zMjVopXNm3MFCP2YwjKXwDp1Hu1N6RNvPBE6OUGj69BdhcK4YUoDf
3sCUqPPbXZXvgY1L8tuHg+nxsnUOW+HsoIhovcI+zhOc8Yz0/rPDaHuClcK06wMvKh6tgtrR5WG8
Ers6rhtprhk94MCjsij/idTV/w742O60V/flC/t5vN8lAgWyPJWoMkECeeFqSvfXzYtiaWi5i+az
vBEJ0LUhBwvAaIjlPXZJzIWVFRvA42dly7Pt9LXVA1en0cUux3EvH+V6P1QgbGMA3G4tluVFIFti
cGEV+6v8k23BoLfisWv9vFBNtun/2sp+IlxciiJjVUAA/fUTdDzfhVG3CoFIhXQofe6ygGftKtSb
lpDYMbcYaeTAEXfgbr1vZuh6MF8eacOyK3Dln11NV3I5g5U7ClLKYr5Q/dILvR53J8iY2Z5XlbD1
yDZ3G47FERdhx+yg2rlfjiEpfSf1ftuIZWs81K/QoTBnGX1vW9nHQJNt+bVan7C/9hivN2qb0t3Q
6I++g0fXAA21bHZn+UjeQ6LKhP7Jfa7UJrdcFdzU2UtpxXo9jM/OFYxUk2FLZSfu8DR4r0fB+E1X
UZQOeqhknslhQX9yJhZFxdXXpGH/F/RWmox0TjIZbXz8VVFc35P8vAERoD0cJICjR58S/N9MXfZk
6yaJ/CkDqDuNAJnMAq4NWjLHTVBNla9QIJ1GbEa/sG61JAthKmjEZBAnu2FzjngfriNEwX8LwhPz
Tjo+KBdESzUi0mbQ2ZrWGMd4H4JiSjlQciWwdzkFslIcrrbLFxiyKmexr0TXJzvAKmkEZZaxu7u9
WkoIPTfAYwEkyn3A0IA/jFBmvdaed6M+fXK2EkCOwj7B13iPGUWpRa2yE5WpNJu0pdgcOcsuiQ2u
MPIQX1eWOtG1B13qWJsgvOJTI7i+5kkFMVdJeLVwjRppS2h+Xq8NTNqcpjiaKVuvgbq78qDaNo/3
q2QdFmEu/ShVTKJeKLo3u1YCx7Rncxn7iDZ0Swl3qAxf5xrsTqkofO6NzaLmrKjTuh/NW05/V90+
2NrEeMqW/fL8yQ/KNFqogOcSVOWLXpSMOCrAIc1IzWklp7r8CLHQmHEuC4dmGbPJI/aJs3lTlPQW
dGLRN9tTEPv+rGWOoxZFXJcIQ/+xWFbBkXtoP4iSxZTTyC49abDq9Yg9Kc2j+FD2CqWtFfUFwS4i
AaYqQrYJgf830PdP47YrmelJ0f1jRG4OhdpeVv6LtlWTYly4NLOG5P9HwWiwsZB2dUCPGwYLI9TY
WggjU6PuQJiRwSCehLM0ly0VgY205QwQOkqD/Ki29g6tOc5qoPLRWeNHoyWSuSqkFuku8jAbf0oi
et8qutN1M3b+dtImgH34fkLXGM+zLYf9NxSwX3fwTh/fGYwNVOYILgPGNT0pPtt+gxiZuYArX7gh
pikkdIbJsfIysFWcoiumBwp5vKcbodzV5vDlAh5RcGWm11jyCkLmoO89x5v0Cde8Ti9K2oS3dg6T
OHP7ikjg4vTNibSr2m7e15CPgUPWJWH72ktAEX6L25A0iNm8GpUPZhnGuNighdy2Z1yXaM6sE6R0
gAnfEjXVcSULdyj6vR/0MO3vqxDnxu7zh7Si45jENiPoGM1vp6+Cn6ZhJPBXTTTGgqZjAiFs8sU6
9dTHxfiKXCz+wN2Nxa/ZRXSjuI2iAI+3EC2XlzFGE9saihf/7Ud+w6xmXCwCK264+U2917SR5TKb
0NfB3FRMbVXVQ1CN2N89pnsQhYzUZK7PIlWUu3ufQOdbk9RMqwCx6WFOk/YkGba3zioKhwIyU4mV
S3FFkJZmU7wPKZ5yjW5URLl6H+xtkCaYwqjPPkJJtwwP8mO4BiRP4fCegIP8AJGup7XTZmnFZKB/
92dis4wInJZhas/V6VWVe6nSj+zexU0wM9j2hBIF8rgzdYkK9Yv8J+Z0thh56F6vKCcL3wRX3MfC
ONQW8MiLK3oNYnF95eDXqiz7BVpvoa8+GkUOgnk/gYPFdhiLhaVMGrcH6QYShwFkLO/9hPbyGS13
vHfiVnDOWYSA0O6eABT62CHbU/i1sLpUIiWjbf+0ra9NSZCYiOYwThYYFguG1dKggrAz+iQ8CxQB
bYw71TFZ0uGhwkM1vQ/PXlwyVg61Ax8frOOPPu/fVTcL4TP3kjQEHYpotD0ZgUCRPUdtardB12Pe
3NoIu9xRfPWbkmFDtZ8YhCbfKQ8f5LAG/jryDgm7PyQtS8QNBlSjy+8Kai/M41ClKgSlUamMr/Zr
L1TLvRSC8iaS+fFjzIVv6NJ7SQxfywerEGMZMyFwc4NmyqezawzOJd3KJyFwcTh74QeS3c5+y22M
OVAMBrAaPLiDolkMHzBTvhWqAcc1Umo2UrwytXclFst3EDve6kKHy48xGiXL8awJdg7rjxf7hfL5
YTE4m/DSnjx1s7OzPlpcIfudZ3HLQvzjUR68OH43Lg/8yCqQ/an7Qw8ZEvWrIOz3RaREWvQBuXEs
YXxJZSeFztSlMmhgzOsDcVAk4GEte8DrFYY/jnDJf6ovEMywNZgB1WXiBUxZUl3YWFnkTK0kJs1w
fSvJ8lFX8TdFs+XrlFhR8aYXIzqq24uVhyeDJ4mizMh5+XtsiE0dtDp+w7oiJ9Wn7DynxeR8LNqS
ZXia9b7H1hAEvXA7WPKLd3ARAHcce43kh4meihjk4CP0edLkM3udqiSar0r+ByS6Vyo65fRhmaXx
B+Md1jpUNIlA32qUmHAUh1kxvDfZcWu+PQ6clQ25ikq84kpBTn5+yCNZEn+WLvdz4QlMpT40F/gq
VLx4pHJPjw557B6PdsisSzOiOnnmk24gAN3G3cNHkCrJ9e9G8zDqHNWQv4JV93JDeS89aL8utWjv
cWcRfoEYzGfWriiWbZBaDpe2jF9TBZT9felJVu2CAfiLok46WDJi1uPEEIfvA90ncGm1WrkFqCDU
VZ5VbNwoHscDovQ9G+nvVTKqXg66zszgFXz7HIgKmi6ycvFT1Ae1sjtVNq4pOwSU+4kJF1IeEL8X
BJfEdZtPU2bFeHi38M+Cbp1XSBATwc50EuOHD90Sm3MTk9vrlHtUrlMjNopD8NM/TfBIeSYHZMX2
G/ebxQ3YnnMsryj2FOlxlpcmFixZdY+n/T8Z0tqfrAZqIDRTECQbsoFOtgIymT8u3eW7GtSx/+sJ
AIhrlhSJ7Vk4Sw3heVyukpXlEOw27D73asOB5w0cauzJthwz6xEHNtcQQSx6swkoEaWsFB7uNi9G
ZrTaQjLMj88t3PYm3rYTxsNrdDMZNa8RS4p0nqHhaO2RPa4GwS6az2BOvoflm5guqSEFfgNejOQV
5VbWyhzgJ1ymT0hdhRo2sG4fpQbdi4n1igT+8rzh/eh1+/3e92r8hrKAMIc/6n7+uXlHluAdrB8+
KkCH8NIVwC9iEUM3WpK0UAGSnxy+GCLCK53YYufOId05FGgObxCGjKQP5XuFF67Ta2qsUvrATOgh
UsO7lv/HUciuN/kp2ETv6mL4d1vyD/zsLojWSBiPPiRtj/0WUKoPxKLbAtlTNm0mrBwsYtAALyGZ
sKQBFyUInFN1pQCmNAL1E38dLTyHXG30pCBlrVvTPf3gP4gm6C11CceAjfHo7jripPJ0pTa7Xftt
SkuVDPh2/fpboF4r/geLSD6cULAkE064KZqjEf5pE7zPcm6L2lx7huzKIr+JML70r/QEulnJvPhv
ztaF1vzqCEv+ipeYKTlIMRGqcwL6QdjqChmLZnDc1Dp2EwnCjV5zmH4jYqe9Ase+MN2cyW4MpQ5E
ohqCr9nbbKpoyRD8uymueEk7a7fQ3ZKYMgTqyjisPwBH+2Y/T0lxuuGRfDSFsHEeA7H/elKstOHj
hclOG60C2OrVNLgD4rrpNE8jNEFm4cI7M0qE6Q0swT7xI4c71jK8All7e+HvY5Yk6pe55AgoO99P
gr3b1Lp/B6fDUTxO/2QNkiwPtSZle/5dJVUq6tnOpHJYyzpH7MW7S16rtNjv8oQhC+k5DSQFumDg
04isDnN4MuFlm5r69qoYGSqm8d6seN6nAnfuu/0Skl6C15/1+eZYHeIMFkyMsNrGRtaXvRyRXDEt
GwYWaefNNAqYRe2y0D8lA1uq0/ruLZ+IknQlMDnjyqNby8l3M+m+jmA9U0QoOwqy4Gbz+3fOjY/1
DpcJj0ARol/vz6R2wumgck5VZSxDEPs5/XsXXc2LuS6T9V6FC7E9MZQERR8gE2srJfV+tgV+fA8U
mN8HdcyFkBmKPfa/9UaGiiJaPknALhSstDak/LTk+lBteC5gmGtZOCyLZ+f4HjhZ9mOFbY9JKKc2
GXmZhgKKKrgmmHB6nv8m709hYuZVy6f8T9KzGAD77bReuvEWGgiPqSpHKw63RQpTbxTXZj64163f
eUD8ANZKOqNDkU61Y45G/TCBlmGXmOoc0lyJs0u5rNyURJ2nUzYvkbUTk5jPmmVOCfxmf2pUQrcm
5PG9FspoavjyvPWGA6uGMiHix3Zd8tQHPQZmBrmCS8TiA1MgewIKYzqV0+XynguoYW25VDH27gyB
SsACxpPu4IBp49d27+s25aWq3e4tbMMiqeuSm9cjcoNcbJFGkza4p06sIYSxQdnTg+XbuPUqM6IO
OvBD/kDPHRiffVqAtARupI4AVY2JfN5TOW3NGegaM4pZ9SlXUd5x0efoSLv31htGfiHLjHb7ql5r
PNqMfR66RKuFWDWy4rF+H4+XlHUrDyn3EN4y/zKJ36hsSl0f8r6zfs0bKLxC+I/t2mC6uheSo0FY
nWFp8H5KA5ANf4mVsRyJ619Is9P+3Q7D6KVQz+aYYh8qts4AGuAKiQPL8jJuwM+LBQ0SzVPzNPrV
u15KK6hZBxzx6Qs+kJgJXp4Pcv8kU8IrAJXIKUuuJJzOaCIdvVESh5t1aAhayu50dPKHTBxtzs+f
hy9zvtghL9LFcjshn3R0Lyn3Q/5kIxAQdSVUOSvRqBIL2hk+yc3vH2DkyXtge5kzqvXYIo5NhtYa
f4EBHi2+H3iEbGafyvS5SJYzE2uvIJBjXA+ovgbIBigxsQ+1FxD7Rq98we7m3e/FU8RAp3+kny8t
bh5zAqXUO67svilmj/FlBI8NZShQz/TeqcNjFcXZJVXUr50gisj3VYe9T2uA8EgptE8bFFf0sm6f
sK8vM1/8PSN8v/p8bhXF9z+z5d9y55Ai0wfnM6wu+mpFo0Pd2zF4WP1uJacOwoURLS3hmd8vcD+c
sKMr245Va2SFiF2OAwvtu4K9wc2LWYEhZSd6asKCOxYbT9Cy4Zej6ae6LPcpi4CV008txHq7E5ah
ZQt5qFyHXEK7uS++o8tucj65e+2p26v/DwpiRnpGLcucvEeuXyMHIiQ3l8nBIkyq/RPFWg43RNgl
z235QWXBRsZkEkZL25zngbZ0Id2CB6faNGyU5M+E8YJtE6kRgdzFeUqsYz20If/CHRgZmgpmj5t4
4yZabtFaFo8KSDcJLZ9J3mP3tZfvj6lUbPwP5lc+PLAnHCis9zgbN/OVQusq2o7nOXHziP+6C3/Y
kk2fapPEf5cRbZCSmimhWiqKJ9L0AHqoRyaJI6KJIc2Vw6Gg7aO8W78FErtjd4B87wUT4DxGUcOI
C3yUwopSt51IVIk95VHQal+fwO+ROn/PEe2MZ9XqegN/Yg4CzFSLmWOAMS8lRsxQyfhZ232MczUU
LCad4S50ejPtNR3aEOs1/5bh20BP+crK9RaXawwfEJNnKM3nA5HLO0DZGW52HjYcA0CvI0UEP/c+
KV13DpOsjuh+4AqthnsULscHTsDiBOjtmlVs+/PRzyFmWy3zClLN68fZKdcGxUaEElFvGc3XwFUa
KKMlN+girZ8tRlod6ZJzzFGiw2DyBFQGMoWFxY4IfjZdBHqJBY3UgOyg8zVAW50oP0v7BtFIpelH
wej7mHcpTJrDxexuJhHZnrWnEcI=
`protect end_protected
