`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
Uvl61+F2jvFGPGXL9WiWhcWb4LzbhwN+9DvDzd4rkxMe5sXaN+2YqDLzFwzB6vfiLUxXH693X6eB
Xw9FFPM1iA==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
BeTt/KsmuO7XXvcPPGcvJJiQH1hDvudia/H3fXSfmZqGxHq5FH69lX6HCQK0lKxlipo8vRGlq3gb
BeDM4WgBEU3EVPMfluCKT/277shLx64kW1YAg5A/ZL0xuFbUKF/8dSZRl0vWcHnnAV1tZyjUWQHW
QvVSCt6ae9p4fTeo0w4=

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
ZJEtzAnBsQJb6m+rRnrtp017n+edqSkKT7Njs3vIqQsPAXEtfVKPZTdMBYBGildQ4yBZP1gHaYl4
HhPEEgSmokGak/A8PV2gLy6DsIJAKXvFMiifZbivOMIXRF04sBnGM/GkdENF9S+jbL77D6Luyk83
w5cWTgAOOUBXMPVi6lU=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
wkq0D4n81d8ZVuh/vPN08pClpOQRlLT+U5FzDOSKM5llc8hH5se66RgXkOQcFk5xPG3+ftPfmuNz
BpRGyIFvvLIt0eyXsuCHTYgJjxgoaLgq4eHPX+o6y1dMo9SJ+LCWChx8a1AOO4l+CMt92cvCcOY3
BZWyG/dm8LsmOWosLmtOh/IpbyKpYiDjrdCMLbiKYr2pb50t+SsJ18r6ny6PgnCHrfqXe7BfsJcL
YfofPZBsIeoTYV6crQeX+r+7hO7QWd2/mQiRRMD2kzSHDG7lGx884zwv9HV118hRRtFFI+5qD17d
7mY6AtYtF9gISAARzMc7bMoKkhD7fiVuXCjFGQ==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
d4l+AKOVa7f+qX7Yw1IpZT2kjhG08YXuNTqjA9DNQkDDpqYPxmpNKcBhP/d1yjBQuVQAqsCwAtAh
eRObpb9GFV1Z8Z7DwUb56x3qu9pLRA0WYGmpvuhbObD1hCUYj1PlSO+4gpkFuqkamSlJRAnjJVUL
BtK+P0Ddo45S+XnIXTcO6IuS6WwDkKfnfCt1qBRmvXpbETKgTC0iRuFXdCK1RXdRgVVO00HNGORg
K/wDRBptqRzxkhKPGM9xj0hAzOnLgJXXTw9gnephIMPJstdScm0ylJ330rfvAORCPl5qVNZHuzX7
QcPqtyGbMIZMGn28GS2YBAj0pGKlp+kNke85hw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Hmj4LHRUoxj0jCOnh1N8gGuBwiXpxvNiRmGLQJIepX8XFpiqMhyFlwLup+O+ovFJYPrq1LMUSAqt
6TjUIuIBD9XZFQ72hVab+PE/cYVOAyej1xneX2sKJG70/9sO6yVvnJ9rzzlEOGjehchm7rgyZbw2
CRJ7u3ZRjIjZQSgb02p/g0oogghB7dfRASzg6BNoCo2T79or5C2ncLg7eeq+dEbZHowCQDP/b6oy
ZoKcxcVNGpt6kfIIl16ueybdxpu6lQ+qUGn2FzXFeawfn/z82bG3nBnQcJt09EWyhH04qJZAe7BJ
HFsybNiIIaXrJzz0aDmEs1nT6LfWnc9bQhMGVA==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 102192)
`protect data_block
HXDL1u8G0m31GTvikUJiEGzfKeMVUnRIksaDTN4bgF1H3h8S0NlBP1yrAijMlkV/2Zcw7ebd0iSD
ilGx/hp9T7P7Ii8ZODFk1H0aWx48acvy0sy6ELXcQDGC1RJyMwZAKY4e912W4W7WZGJp+BWjn65j
tejsFKDUZTY8E2Hjm0BtelqMF95+YCD6B4b3pBL9TTomQlb36WcUe4JDHfE+YUcPHUmwFSFt+jMJ
+L7KsV/WRZteAn52TyQTl6r7osjzPBv6ooYRfUXkvQ2kqrV1gAA+ZAMDFqENvL+l70YGi8/FQIac
tm7d+hKexx+Onj5cp0oGCuEh9Bv6+JMIfONX7CYHJ5Ft8AW5i727DetvifA/aK5FQNV6QZrivbuy
0S+uNPRVO/SsGMGbxH7v4rwe8uim/sLUYiZSbCVlW6TOVH1uAf1FofHiDzYgU/xE9QBP14378zSH
GZ7yvjPj7+rjJ8DKrpJnG3jwFkItBpqRPDhb7MifzumvsJOKoEWiXDw3lDVxGNHdE7dR8skZxy7K
N3tA3BAJjSdXNRcsQEaASo4LGPoXxsq80h12aYSVtS+PJaMm8DZBLaJ0PpTEI3F5yne+IRvb/KvS
YCfpRlW3tgjcvzgQTvJ8AHsG8uEeh7VnCCg5/XuGXdxvG07I1zlPW2fT/iLvEFaZrFBRglmuXx5D
z7SubWVA6HKWgOQIg6u1/KuO1q6WpA7s7/S6enKyfL7dIetnbrGLIF2KPMQW+pUfZfF6n70/+Z8q
2nmUFh/RR5G/4FNxEZEyWMcUtpNd2mwhBdPANPpYVocf3sJmk9hdwL7fItSJTiKWY1PHDRSeV6dP
vaYY+ABwesEvLuNxNA+Y/fYJLxaMI1uMnV6JD/fQVW3mtValCsqIH4acehr0ZbfKvoux0sKyAo+X
AH2iR1RM6Jp3yvW3qa9iX4XDLkaXXo6p5bnStNbtXBxzdHwRObJtz+AxmTdsICS0jMz7w7Dr39uX
z8LCag57W7A7MDv3eHj1oUcfdbnxpoCKLMYXlirbRicsKQJ6sKktnQlJjSCQWDRoLiqq4az2PmC6
8VqYfoCGTxW5J4k+wAxU9VJxq0vKqxhF0GV8/e500Ay67sP2MiDOp0TBrz/9oG7P2odVdCsjhscn
vLCiW7mdQ3j22r99/LqZoT+VUOs0pyPjQ7Qm1Xtt+aYh3bzKCxWBGdoW0au3O8mA+LuKTGfH6d+Q
mZmuToOMj2ijE7w+Kgw/mHdsxDoHBsycdkZJuFOFQ703VjxmdrX/F0z7x/ki88Tt/4yWyg4w89C2
BrQGhGhHzDtcAubv6qCOUodHZ0n1J1LzRGcrRHso+gM+iY32t5E627DFNt78CNzCXbwryIDnuyoU
ZJ9cS5lFwuBLWUVnmS/mbihBnPmF9EZdvmZJkWy+FJzpvFAxq5nxgF5Hx3RzZUnpoYcFgu04fozI
GgcSvxRtu3o4Dw9w/benjbDUdpow5LZWOJcZJq686Xvcjf3OhniQfkh3CBrCZg+EO2mFKLW5xVAQ
sg0xSB2M2do6ydCNTaUopYwBwLR8JJ+Isof/TduRfIeW39N831nlKmEp0sMOpEu0LmMcrC46sgZJ
C/0UMOBkchX1G1gj0pd+uC1J2a90s6E2aZhR3H9ZKclUyXwd/UHrbJgsVPDidZc3eZ27La6z2HaX
FahA2ODzAqjrSOS09W0TKEOdms1P1dR4+r1QGpV9CWKEkKG8H8XsgwGRsC/aK3XdbFfsKJgurD7S
BPSCLBw3AupP4k0Q/4jQA8Ts2OgWtXLPi0Y1CH4BRZ8vc3KX1xcc45/+XsGI42L9ZWelkbgtuvAJ
Du9J86CdzdTfXqJ0gbcevcNekp+k2hGZjmWU96Vz1PUjX7/VG5TTIX9rNSq+Rk2FlfX8+77+vGGQ
QQ5e+L1jrh3pzou/WfwFM0gFGKOabqtvIjoaiWJHHsuXaH9onv+HbMR1HpzN8/6n4fwiEKpPXGw6
Im4q4eZOi6lwsOhfdk/XhZ3Ok9YT90RLzTFSIhJL/tgNPHJXc0wXHoUeakqjktd8Nq1dB/b8RhiB
sGbe9yWCdnFr9Af/XzBGvWY0LArFrczXKirGlAmqKcCjkgtPkTXWylLIslKbE05g/7GubDh8TdOw
a07s0YjGSdyZf9yPlO8rsmQ1jPdtIxpAXLqTGtxu1ZZfK1gnH5qykyt7HmzbnS6oGqmf+grFZsoZ
pC2BK7mqckJIQHZwbZgTv0vBMxLzu06PsDuzA+RvhBWxlT29Avf4A/hzqckaLSrAyB+5WWWHjfGy
qOPrxcABocI1YCoiTSdu3ZlQxJZbDXHwbUtSM0gU5D9rTclXzP8W+PRFVdawraJV00Czticwr1ll
gHVI/WhY5cYs8LBiPYZCIGoDtm7bNlSFe79Qa1pdOYsAxVMJ0bI9WdOvAfo+77bfS8pGroeT1YHq
O4eJ2epG9Gqkx1KqFIu1iTA6mlieMCXinUadNdGeME/lO+y8a0rCZOuuOvJZugsG11X2HfzEybGS
/AutPKdjPKWL13ein1iOzCYxJctSLzIadAUrMsPnNzqaiCua3zdxNLiNxrX7TwKa2kPNEZq4/T5n
poNoCdlHVoidr5erGaAzTpuA6qhRRUvPqnw29ZyB5PufO15l8hmZHYwJ5WjqX9UM6Z38zKJm3kGv
L1hUHQmjCpVwzllI9V1KQ4bpAMi9OEJ7Vd/VXHdGrR2WqY+ht71kSbYqxJLjF8bjgrQ4UxBBieRH
37NGWxPuhJbufRHjy+x1oXJe6jFxI0WFnodLahZrvcHj0hWx0GicRRELGe0RRy7KqtgpUdPholYZ
7FvkTLLwNy8lYYrKKGeid5nYQC/uetufgVSFf2t1vUrbm+4rS65ffdD7Iq1trqfhsgJ4FsdJzbhj
zieN4a4OGQEu6BoUG6Xf6aa8I3k6QEmB6JetqzVZWy9HCd01lDnctu9kLyBf7ZQimWZ+f7B5Leus
cTtIqdNk7avDYKAv9w/vvVIS27x1RqCL+2yaW6S8Dr86VYc9TfdccrKFK29slseM7/jvMS+V4L/v
K9QG2z0lD+2QuTvD8MOhx+chWg5bnqFnrQOyXqELXAUDyB4eAYkkG6ycclxqd/juC83U63ZYyqnM
AJT0MLq56QC92PSc5q1Xbt8R8e3tXW822cjGNmeQ1FF9aAMbNxorEh2wj4uc7X/na0wnIh/exn8+
spoyTx58050GgSASO21bwKOV7bfiFzRSIJinb5uGyx9nw80YFcHrVxgbuh7UK0R0QrbjqFT7IBmL
NEnyL5zBTDWWvfq8IcQweAgcXIwl8YUmTSTv05SHO3X2otIltTHFSScA67Ff+JrJscbw5sKobbKs
uT5iXnrqKYq9f/U2McrLgR963zF8mf7pOhFGIrJwnGevu5yAqOFAkbh+BkRfr29qfBsPODHeecQs
iuZItp/xoAa7hKWdkEn31rd73xhq+howHxozsMT6r+NPRO+HORz8SSRyyJsGBRJj55Zu5l14jnoP
hkzhOKjgFUZPeDCN4VwYb2mazgGRBwR9tdJKVgZKXanQeRMRh2f3B7pvHgXbTNG5rN3LQdgxDelk
RiFpLP5maG9f+XVuwBZRX0v5ErXU9zMqnSQcBSvdLl2FoAjENhVAepnIIQS/U0M7D61tFLpsF0X2
nYeGkQuSEOKASIQ0PahxZdzGYpYO0+FVoBvDQGMZErquqjsxF72Qn0k3uN7Md2+3fhJ0k7okoEpq
NsRySTn3wyyeYNRynqfO5tFwAnoKoWSFvhgeuRFgktk3dTBJDaHNWoIg8NmVDpCZ7Zcnsf7BdQYM
6dWR/U0ulDBqeaFDoCxfWdQEY9tialUIExYYp+JTn8Q9a8x8Z9CMoih3m7ZQPqB8eW+sSobCORDb
GbWzVWNek8VPHLwJxptM8mniV+nXZSgUmF5dC2jb3eu+C9kqObNGQA7H7ufx7hzyNGUM/phkxdLN
u01QSfq+7s7qI5jG6muusPcWpmNettvIjBaE1z2Wd25HAGkio+loocNVHlvI0jEgiEVRcrq+177K
FyWhba7s84QOY3oaVCFmiP1lerv3E6w5CNTY+I823VbEGBwivpmE5HUjLToQv/7SsDaXjlQjuEJk
f3mk75vuDKYWrp7FxcCQWFyG/QA/MxMHhIPdasjV177JleRiiuEwpRwdRQ7lEZk7Ihd48Td8iGI9
U41XvSXbVS+cSX1FvQ0dqRIwTcxcrB35npV0W3ebNEkRvoHoGw20NP4e2hr8iiXmrx/M/67sB2F+
FkRV+h+ERsChqnvbdR5HdUbuMdc5eYpNRJiFw1VsmqLbysSy0dARSsozHWNNgJJ2ZLhU1XRISfA8
QEztI3jjjUofRzTspkgr9TFGGTw5YBhD2StG9NzHtKHBaZer8f96YyxY+8GsPo+IiXSW6Bh98uqG
VxZ76eEvKQmvQHnDzKiiuU8Q+35IIOHxKaOrV0xzo6KHF2fqiySaIzGX3REbKwNsLXzXtzw4n5xc
/iBUaGlUgY/SoWULBwAHHif8AcQl+4HVVaiXRdI+02GdYXH9FFIWlTJgQFXrTkBtiyJQqm+98hrs
5vH8kSDZwykm3S8v0QN8lId7RLuMOM+X5kccWo2YCUHLdOgr9SIuVW7hsoaJ+JNLajy9vDWfQqHZ
eXUKv36g6dQH2ja1xn5kjn1IEK9Umz0EijyUgqeRRnT/ze5+xqmM3k3FrSvi30m02Vn9e+f8na24
zEpGELnK2YdEcMjKyOJLRC0DU9z7AVg57tOTpDHMMMlYzWfYHbMqjfp7Dd/aw1RlVKQk5NLyJtvQ
yHi4Y/qDkcXIci9tX0+n4SHmqkgxGrhXG03o5xajMFoZTSXyxbHH4MavDB0JMk3knTMefD8W5BGv
6wfzPDiayZ/P6pZUSWH3hHujO9Urnt8HJWgn4XJDWN9UJYHqEN812U5DrVlB7Wla1RQPN9M6r98J
WdEKYgABJGdxTXUy8ov4TyNK/mJEdqVjQGxw5BgYq+aBn7ZXlzIu7t8zee6lF4U14WdPgzaWoSA1
dN6T5RxUstcVIrVnGpnBLNUQ4RVBkvYs5JoEk5zyIelI0UxdKBINj04rPrC/e72bwO/Y6c2yDDu+
2JaFHQsd54T74klafDTPDK7L0YGWEweakXeu7X+RY3agczF6Zwj0yktC41ylojxlI244oHdUOX7k
tQjpybgaBCjiVY9G5qxPU2lB5NTzHdofT/6WGtznGm2Eh5ff3fwL1YJP8u20AALCKCKpXg5oXbX4
6gzdrm2qcY5Z0H2omGs9mBAfZ1Wlej8KkazE5eBa3ScqNx7KsNyn1Vbre6zo0NSqGo5/mJSkwBmt
/sWsvK4EGofHZSmIEe0hw1EZI2wmB8U93MfbDAsZKtFTCNEZwLdF0G9KTVFbbPhJC0OQm5soA08P
xfWXa4Rs4ZSum7MvBMe7Boo3BuNm4E4H8PQf6zScLpt73kXJqK2KJ6M4skVx/HjIzb2KkHrlKceg
vQzctZYt9FB1FbEzmU3jggbqOBnsz3ofe2054x1OYBOlG2lT0qiQLd9j3VUn24SsDM3mtkhzmOLF
lMRraX4vXQp0u1iwLmERHp73olOUFjqwYrSkrgKKXdhesH5os5kMTon0pThLg1NjhG+JzZmvgAMX
u6Xr+WACZN9vcIEJg9yd4fR+lbYPP4615dYeGe7y+b7wVd91aV4OTL5Ne4ZZW/Hvvdh5LDKObGOk
XaS5qFgMPEyt0yknkHxtcMt8ZUqi4YGsDoHX/Cqb/p80ZzVTQ4/hDNNkymygr6yad+IyN9nDRiWz
Tp5n3EmykVGVYgCvXlt2DlOVBYmf2puu9tF/YIiDeSTCFPOJBdx6ruYmunThlwsTuwWPflcxWhhL
bZmBI2m6AqDeiWaAwTEKOChAuqi7EnMXwhfVIaRwO6ad4ksC4lqI0lFTik8f/fWIFybVp/npuElv
MEdckvQoExU0pbUzff4iswJW396kGHTM31PrVzk4rDiCw5+hA8OPP7TvYFe/Z8Zu9PTfbwjsW5S9
cq6vWLpGyKewt1ef7wy9+/4BVDY6kbG0R3+OqfdbCQXhGb8rC8y47Le43J9BhJFHZXZBz4xLG9RQ
Zf08Zduc9HxzYiWYr97BdCymmje9Aa6rGmTiSsUicqk64N7Xc3lIu0Ea1Qpu43KOSwSF9Ded4OQA
JMsbK1duyBOr4ZubOaVSGweqZ8NGopzS5NrWZKILtfsb94liCipk7vl9i2ucQj7u521Qi39qHTB/
WLZ2jh3r+msLDGlkllH+zFlUny8kR7zYfPXROPAJUNJ+4HGiDEN6L08+rAiS612+ZiOMsXiCgEeL
iFIRRa9uP0AtFHeGGez9T8Vog/vEGJlhl+iJTDLcslt60sffiD3WwICcUDjNmDuNQRslyTVHqskC
A8J0DCHPF2vAyiAVUS/BBBlpKxQ+h7ONPHMeJ51jrdWlusO3bX6dFsemLs5tuiPLjqxTl58+CZv6
jgyK2zrHWNrzxwDllVxPCeNtC0LeJLtWd47/M5h181gkj/EtIgl1UGJNTrvhnlacxFMvRnb2JA5U
snYDwNUwsKM1HkqtXYVqqA0vCBzJvVRvG5dnLZMRK37Iw4cInNGiKJvXe5aTPZNb1qQZB0Ri9BVr
NS4oxD3kU0S88ChkYhGT5M2xrzT/KgjSJRis5tV5dUsDhxm1T+a4LOSSSimKBzgLSYskg19C0XH5
6C7P9N+rSRGuFtVbK/uNIE/v7b5Y3LbEUOb+KZCJnwvErfV5PXblQPUi0A96HGfLGIjUAy0gseyn
cEwOUJyl1MNszMCtGSnug7XyREVd/jAhiJbsu7Acc0Fs087mztobT37fDa/YMGHEaBBjnTeJdQK9
mlfbUhBu5KT+QVyfzkEnVfR8gtoL5Tr4Xea2DJyKJsA7z2LTEt9Zwvp5ZXAC00cW5WAJxyTwzOWy
Ph0VhZuwmkQPF/mYxq9Qkl0Ym3D4w9Dvj+rlgYKsnxGwSa3oHHZmRlF8onty/azPPRoLZSxOUYjx
hr9fPAXBVmA8L3YUmo/IbEQgU8BNYPxZjzrz0LTif8J/dHDuiEdv0mAED2IEUEJqlIrLChIxtj15
/a6QvTxdSNqEwcTSU0chgIN6ONg6BPiNdXREEm7uzToA8nCSzj4RHscxcf1vDfJyhGihyNzjCK8+
lx5WqBMt7V8aaPaRVWxViW5SVjAONVGDpDiZKyQ3UerGHIOt5dFFdJuzAGexCL1PYyj8bH7OcGeJ
cvo0cBcI8L9u1bMVhfLkIrc8vNrV3jvy+9+AuZ8UsZhoX7xOUujLOgwlSbIlFeVeV3NwoZvbeCqi
p3N37nwZjny45TiiYVOKerK7B6095SX1btMog2itKVNUidYS/nYj4PC1mx6U+aCJlYr2SpQNGDZ/
z9QIlXAcFwxczJkf/xKIYHUcfXOPv9sO74PffSgchqUdo0vbi7x4L+cq5LVANyd2uar4KOFah9Uz
FBickP8fVb79wqiM7SZRdRFsZmJvA4XeJFOdhSPYUhcUFDIGOOYUpX30sm5neOwLV4IaeESu19Qz
yirxwLk7PLeI2xbkkoVFHYM7uiHjKZq9dWcwGCmhz4XECoMWUKsSHJIE0N68vINRhR39uqq/Ldup
I+H5/m6JQts41c+QZdQCLXmTRYsPZTxPh8XRfApomChOO4KvOR8oKk/F/ZYdpRkeUrcEel+oJJLV
TXmcSJJAwkoLxzrEl7sRnnBu2fBmaac3sO8AWJw9UbZQM8Gk/suv7PpxuVboS9ZtEgSM+4lDaQzX
aMmrLiL7u4oJBQ64o7aTh2+tt1imDPil6hIUoWug4NLFR1/3ZY8I188QILk6mcInVQPc+WahWcPa
yXNVu9AThwx6nu8Tut+5z2GhfHZZZtIagQXoH+w1ibuxUs75siqnErxwFoThhyTAMtI3i6HqzyrE
zMrpMNULMbK97xHty+7vXtchkWP8TT3jw0nnxrVFP/sOpSYfaIFeXU3gvvWbXcqAhQ3a6XaTiaLZ
OLbGFad/TE5hnk1pSDyIEZjW+mdE30gKZNoq9OUC7w2wYjD5fLRBQdJMq5DZ5SESqq2i29rm6Px3
6smXOJsmEkmHePnx5DO7muN2SBorv3EAUm4nlMyMmKEnXUk2MYts0ylyw1mNeLUOACoFeevnqXSU
dhUWuV5t0T4sgIiyKM9nANkrY2Oe9f/dZkcjv3/wKNPiA4tjsK25/PkUO37qcM9+wrhfkI1pinuI
9++7celagFFpKyw53Wn99ugkcdK+7f85SOGlToQ1yEDPQ7mi1bOOIDZZNmPSWufPauS+hYzf5NGr
QPqOS3jVAthuTxHRdewR7JBSsalzRIG+FMOBYB0xBI4eVkO7hNigAZBkoPtH5XPWWgQk1d5MvQeV
nl4JV0I3n6EgwmXE8x+nhViOOjxr41kd7dguNhT75lXcg40YksIrvd1P/w4r2yaxtNYXVBX6Uadv
bV2ZhduQ3ODuswn53qtFUqhDOUKe1zJKXpvUnf9fP0GEvdg9d32xXmWqWGFCaNK3ZBiI31RLlS1W
3MQF3udbvR/PtSNsQ7lyXiCoMxPnRRxiPHcjLLTnN6iW4JeGnzZzhMfWG/uJxhirRMQT7TknhRrr
Jto998GYyXc1a2bD8Hpd+gMyxBoIw95t1RpE9PsjYipD9zbggzRWu3n4K1VTQe3FGfn1p4Sa6JLW
7TG8n6nHU+LKHx0+mgH/htNpuRd9b2aSzU5agoTq6XKnkiVafPxitYZQNVAmFEuKPlAeJPj0Qmdy
AK9E91ap19bbpvy6SI4GvFL3lg3PAEcFhlnO0c8nleRdoUaXbK2qmNHraWFJq6xGLH5p6AaCICI1
gjquf0ljXSdX7j7kA6fbAXLLth4KGhUiIeEeijIgQvaqE7s4MGQpw6bj9p7/HCnfvlviNxANDOC+
JzT9LOL+Ba7eRaI14GzaczGc07+PGZDwFIpQw3iyTQj6QZxbXn6Kv35Ey02TQq5cSA/sA9Ml/3wu
tWXPGqZEcDYwlCFtduyQxkcc0HidTMzV+hbbCcMxsaElIwiE694EwFGEK8yhLem2oHUX1OYqO9Pv
QILvu5Dc/Ea1vQfjpnA2hKZDsd6bvuozJWvvDh1DGIAjfXarc9tUaFBS4kmZzkou6Zl8AmLX2xXk
XFHUI0MWfz4U8sLIiRrgsSesgI/0mFXDlLLgxel1JWFVzrWBkmeoW+674d+Szdc5msCiEccVeFb1
S+k2wth0jgs+XeNS1h0K4H7vy1AFfGGoJjWaxMZz+VOWzuVj/vwIujjnMvFoKeS0OnedirUCl9q5
XnG5SiFV5DyXS1L2D0fUivEyonSpNlt3EyelIKcURPAhjXimq7f8Ei96HS/G8SmkxQnBAYF6RO3p
Igft5yNCPpDmrDxMOIkncAeyuaTRbKXWCePYx2fNPntZ/pABQUYC0eMZ8DsrHSZ5Y+IsIBT6Rgm3
eoSoJQiCQMko67xBwKzngnGzArRZcE7kguUkVICGNHdPj8xiVl3tmqRgHORKc/qI53aITJLx63nG
+VGU35kSZrhDdoIZoLKrV6VKgPJUhjkONqCE2yWyFsFa31jbuYCkLGVVDev1BWC2xR3RPWbF7PDI
gHLMmd7U507a/W4UWGv19HrPkQnuwee27gAxebMC0zNaekD+iWVS90Ug0ja4wars643d0Ns+2DO7
Qmnx9WLyX8uQAcz8VGuCxtnEnWg1ZGSEoGdoMRduhfszRIcfVSMoDiwCRBb9pe/l9GTCxJLJaF6+
ZccruowHxBH5CsVHKQfG4MrC8hBMqauz4tXmUE+dwbNXaFD84M3wWZ0AWO87hokBkzR9n984T1/U
aPzhdKcoknoMfF4U1xtwuT6lRRMapV7AVV73pd2G0akU+vCTsoy7EtioCUjJH2DFAmWsbdGwKL0P
B06zg9/WSF9UjW+N7YUCAWa0XzCVAK6jDZkHcXOc0A6yb4sFTe6koFOiJkeAk1LIrOf0QNKaDq7g
1uzF5qCEVsaCHr9Vpra1BUskchrdeZt9npCOQNelzjQ/LimH2epPhUViwVLsHHTnZ0iBrS0lzHmF
JYY0P7Y93xHdsTHnfjp3opEozMpW0KFQxQCZL8Ow/Ii9MaXj/aHPl+8fIVLSmVP6TRpyLWhBWZMg
KVz0fcW4sqc6cVqpuEp10skGW3sp1sRtbEtT3ccHd9iPqL9WhCefAiqMeV27q6osaJ+FERQwij8K
npd3SO0KeCTtXjlcsInKVB2hoxbqwNhK8uknIyCZIJaE4fvW3dUmNKfGjPmUOjglwAxhb7qpiTUH
CQtDfXvgAildMJeZr7Wt9QBKW3xtqXwCK42oHznFHQIVwmIh+fZ/yEsv6UE055YkPzW97ikme4yl
ICWL6fbaUdmQBf9iDtoT2IluPvSMqI4g5fgY/3bTfgV8FlqMLMYIMukzgFxUi2P+NQ/DZYKXICxs
Hm83naZtQ0GfU8/PACaa3cNZDxLImBSARaELwipWrEKUjkMhMC7AW9UpFMofb1POvzHXn+qtjh2x
MHfSmbI+1j+50i4zpJllLddcbmP1Y8PhOQrvKnHElXP3LrdUZBAv2S8laoIYU5n2coG2qUi+shgv
S7jctr7oIob0DhcVI+yIIC1HJYV7bcw0lF2yTEK3aoAuERP8dIsRHxJ/fMg9NbHv2xaWhexSdB3g
to1q5NlEr5QGQWHZASqMAR5mJ9n3U02Hm1zBig+MMDMkP/vwiwORJnCsXc78lJdkIVfz9lu6rXVZ
TvRvSM3wlieGJ9JPYk7uaw8RdrWcRfTocZAvMK3CtSu7clfi9fIZ3CSj39XFEboFVNyWx0nRv7ye
HrDZ58w6IVSYm3U9evXCPKSkz9Y6sGld1vUlxRm1NqrSJt2/QT0SBfjHKiu3wgcGmRe/1mLn0XQe
qCXhkMaibWW1LhzkhFPtgmBePNigPhFNYD9SvtEw6Nv9IJFlsOS78V7zYZHCWauGgNEnSmx5z/2l
BgEZ9YXGg0P7veWiNiL9c4H6g3porIH9051uv+5ImkU5Ws4CUvyaTJoJygzekAMzIj0HoT4JZ5wJ
KXWn0JVDB0wUXUwB2VX99KnImbnGtymmvUBDQl9O0/CTJk6kkvbT88v/pwh2gWGP1TicpO9qj1fW
8UAA+cVDti52Bh+qVDBd25RMZrZBtcpdwlJUzJkTVSWqwrsU9xC+CryJbygJKOCWvSsXoSTP6REy
2qEO4RwE43df72l9bOKisgC1lOtJV6E/Uqwe7m6DSka6/1x8Afc1s7EZEpI9mKBJH7oVAUrmqB/C
v1BSCZOcLfPuAvosKxhMJh0jWYtvR3i+oaNWc4mnJubnRFR5L9pBjSDME8Wf4UKAYIgiH9li5bEP
Qc/nBymZOr+RRdD+ft6cIwpOIbMmxW0ckLbwvbqvviK3dvmsERxnG89ZnVDKvnG0MLCq8Dg8hHt+
KW+8Haeb202+tcWZRuI5SnyPntNyfWFS8/GG9/nqUkfzM/bu0M2wfs089nELRd3vX1f6yae7j1f2
RkR4KFPKnuiidgHzNl/dhHwlJVDzY7rgOZEWRDZKC7zfGB5nTYUDr3Axr/b7jM2rDe+SWynvy7OI
zVAw63w77vRPgyDqvZ8QjLV54Ebrgn/1EA9nYvOo/rSJ2IjMc3E1lqmVAMS8eHVSrsF5CD9P0Q8D
rG5w667AVPrklVB/1K1ALb1gEcWQIMdAIGhUOGhx+xUusdXcWh/NyL8/WMLGtAfXAGXtzGD84F1s
f3ACiUjQ+Gh1XU+fPEx+FYNM8h32AF5KaDniR+P1fe3Tegttigs73i6kPCq8opnJbCaD7Rc/RdSG
/w5HQLTnIY9ximwzLLpE4VFI8Lt+V8e4d5wYDd7a22ioUVrjrNOeuyVN0QgKRkjLWnasoVCyPEkc
P6HtqeDRI0ERtfaXGeVltwOxsaKLHQQ1EgkH36hkDvMXRFYgWDPOr6lzBlmqTtPK7PJg+skAHv5Y
oSQIVG1hQoe4JqVtqWPBk2cUEE40+5seOi5KQjvhZHvijiLM5kuj5QKtdJbjpbgKFfkqySk0pJp4
th0TK9X9p3WqXxwQpbcies6bOHIy/ccFPR86IB0Yz7H3bXMR0aUsz8YgcjUT4CKPaFjEvs736Njb
dK9ABJ04tSHebW2XugjkpsMMfivRiYpIjmcBur809WUUVjlSkP0pArD8tSpfN71gP7buy1YLAfTz
Bgkh7zko/fYIt+O4ICUt+MAJlDG80XpJRQIfGUDWXY56pMz2g1nKdGouLM+Om392Mzq9bKgAPfVh
+dPG8pwF+Ll0RiQ+EDVhPtMvj0UyPj2tua/N1OxgHvNYHztwYSX65ExYbQCijZ9aAV4kF80OsD59
AJ6/ZfYeKtGlqeaDoRwBh8xDn1hWspU3y+pCJJHrKhQI19iQqxmRrCoVfZUNjY5stlOWNsJFG+i9
oa+f9AUd7Xcd5zK2KFet/vdfHugIQHrQUutzvAiZRxYLuNTUpxmGHxZNkxuk9h8ve6PuSkhjzGJU
SvoaDZLcZIOHTcgO7/8/+KK0/Ml853T2V8GltbeN6EBHTdvlq9hayT/m7b/dwCqFmuvG6ijz7lQO
HAJdcJpi3QcW2uJJTLIyZOCS2icnOXSsr0rGOGJ/8+8u9iHDyL+sc9TMt4ZylCOE4YweAyzESNRj
csM6Y6S11iV6gKQ+2wxP1IykxAOUUQ1837RrjZe2eXuGiEHihgbN9WDp6OGsyBniePyRArLUYWj4
xhszYTB/nsQuLI/JgI16LHQfrfkobhkD747wwYuv6U5kGspGpiD8yCionRkaFiAq28fZYhjgqs50
+3rAfs+btuu93zKO5rVxDpq5MOfX1AAIWFYzUJUpZyj8LB6Q5lpECfCA2BMRIuMn3sLWDqI/HdO7
OAJL1PPV/a17/78zBd919yo+JAoKyrpUe0KwoE5q9K91dDJl/DI4NzKihqK0KQDea9OKqjqTk8et
PtIJKGit39pkMnCsEo9HeOOQvaqZMI189mPtiyg+spgONhdWn9QZQOeh+j/ad377P7fXtLA4P6so
PZJHttIjfeWsMHRlp4BR9uDA1Jkmn0D/d6DpxEGpGrWpvFxtF/8xLe/xRTKW8GLX2fDNunhwWt7L
JlZeBTT3m6D8xZnOv/DB95WKZ/EicBioMkP0lDCxXqcmFZkwAnJT2GIMyFmQZZ94J6HUaQs60VXO
VXtRtGoXEvhr3m+Lz+6PYNy+q3LnqN83T4UHoGxoKoendtS+88LmJ/zpmuPv7aSE7QtosMoblk7Y
SU16tPGxxvWSHMgA59Ba3/fjKtoPBEK+XohBQEX+uieCIb/AT2nJhsP9VVipj2BmDgx5+tMyHqUu
Q6s1WaoEuLy1AWCjjnV1Xkl6t4ilqyGcdEk6rHXiqYbBGHIMPCzpXkG7bYouF/27WM+aHvnIlauQ
TcuhabGHPiKT9XdqWfzYCfxkGiAI26468sJQIx9x9hZDQqi0AbhWV9IZB3DimV+oT8vRnIUJ49SU
xB3F60sLlwQdyaggZGDELA37IILZzJfr61q3m6QJ1MfRva3FlfDOLHWSqmX4mBFS1lLoJHopwolp
obHJeiJ/PFPamstUWAtmWptSw8Xm1ARxu9DJa+DZVgKLJ1OMhX3l9x+DNhMdt39Ikj82XEYHud1p
oAfK0vfpwsBStyE1Iw6D2KCaESMphwlYERxl3o3P8+scAgjQHdug3gDgxKvLsSN9OunM9Y/kBnJ0
/7hL9esRD8t/FKdsLioVEED8pjfWRCN5cViNhu9sdzp6WHeqOCKwwGsgnAA8IH/hh67N6ZFjqgoT
nDk2FOtFD1xDaWzsotnvMHvyTaQGZYD/REf2EprTJtbHAPqujF0mfIgDzYBY2A6EPL5soaycd4+H
F6yqIgiNNvfGj+YkHILE0qQkihVBAJ6q38H/9ngddY1tM1IYhb2++PrZIOYUlAS1VfVUF1FK56LE
sKg/gRTUipKbwlxLUpZ3gBIi9s22/wjSyv+jp03rO2HDYjVBZwYKgrtsDvEAe3txi4JOVhZvRuPC
cUsOgnN3lr5Z+pYDRFt3pLRErMAGyT7GlCSRjQknr7nSCU3lTKEIp5K4qb/Odlyci9mZbA/mHq5P
ZQ17GTU6Ezvs4zoj7DDGtDuQCpkT8NYejW2xZ8zmPTrpLp66l1zVnsfGII5wAc6J/Xer/utpPwJL
/dfXrRymWOf1XZjZlmdmCr9HODa3EAefR5McXZLSwWzFrIn3cdcevW1mp/VYboyl9I2ahMw0mn2U
DjJ5sgXMy3JFvyUvktut5GXsy3O1NwqFeJgAWikEj1dKEJesSwLvbmK/tt5/GCy7PjPEYFRtMLkJ
nuWQE9xePfRpO97q+lHCJMaiflDEBfusYuum0TjmLbNqkRs/eajxUIHDTG3eCKhvPB821WLGODwl
2lgDNp3gjSBNe72IlwyMUqhULyNYpGcVr7rJ2bW/teIOVfVmU7xJGlh0oiA9iGluTIKbvPma+pk2
jwiOX/pIaqne884PFg80BXAdPMxZK5fubDgFnX226V5GfsFsQ6c8gexq0cGP52hIy0p2SUNgfDSO
th86/pB5V3w8Vgq4YzEApva0QZB+Gos5ZoV5cwklqzX2f/KcJg65ibDd2cPUdf7/hDdhRqVmj5AY
xbrwrj1dUK5j+eqmHul0IqetRKdlnD/9xsOLW8h3mTz2uQUeqbk2h6othG9kPheqAX0S75G1d6l/
B14O9yU5AwZbv97e70ueanI85M67aUvRkTx3S9RMZuyPv+RRqR84SuA8l6Ae6+uC1PmzqNEsrnPY
TD9fAGuHT5QCxd5KsoBfMvfWkcK5ubUDNuKojpV/YfU1ewu3urzHaXpqWAlqxox/ZbXbi3whKIFm
sJjLU3MOa0YlqmNYO4KHnCDVpEUmN2hl+IdqNpeLFZ6UlvRzM8wXRr44gJLc7qbCEOm1yDgk/ksI
s/MoOB/9S9xhtevpjhKMFIppxAG4wXUaw0AaWXA+WjxlbzRHBqVMXV3WsljUB7RhVRfev437maIb
Mbi8DSrWNtTnTag5MVXAWMmLt08sUMls1tSQvxYICIRBVjJxRZWQkp0S5OQ2wupoDCsqFAet+Fer
8BpS59W9LFwx1ZIoJVxqRPvLqkO8m0bXmW8RHcabiOdRE5pfLlvcFPHcXbvWTnNBf7Hw9J/SYLaS
wyR0fSt7ggdj3fdFFC9a2ldIhypgQgT20cnegAb0iuiDAug8xLdQJ00uoAFEEdME3WjNM8hDNSK0
Xm4kv1GusG8a0wHSx7hijzjE8OEeSW8Sf8IAtPdtBjvepv1fJZoC0kNAdP2ouBm8SUzT2NprV3aN
Gh8X3Wvp0/+w+4lEG66HZtCpjttbY1nUb/HpjS9MS3KhH5fJyoxuUhv5XfjpVb8HCOiRaRZeMkgA
oyxH/kzbSMRtv0r2ZoheKQFsIu2rGQO4ipCbCRP01jb/mZAmQYA63z7ItAlaVf8cxcDIjaprkfZa
UCBBJ5hTDxPPeMTYAwkjTSKVj3tB2EnaQw8DpPNJcNoo4Kxs1OAhvqM0/BAicRBBpcLy/pGG7Tpq
8CcIVyK2G8OTSbrk2R9gXN6xT8m9EI8kSA+iJd0Qg3fjTqrKVYtdYgkRvYlkH4SivtH4/ITlVvGe
XBqbyzhEnqAGUzH6OekCfIi/++3H1GtGWm1oixhDCWqP2PmXekkiz/G/KlHC1z9Pa2Uvm2KqByJs
aEhztmeRQcnbxrrhhJkCT8V+iQstwwO+EVy2fZKfd8AbB6BjZb2Dm8xtZwaiORsaDEIDA81CO/54
mR8+NnECk6HeX0bxZexoP3HH/v67xSCLgUReWDjGiXkJXrbpvhVjozazQoTZWbuAAFSedBG1bRLJ
lKa6mE/1rHXW2EVRFFV1LJrNmLA9XtgXnopRHry2DJTgtcYZEBPEp5R2AgfPwdCVP4/RlXUXBIDh
po3CJuTPQlEvXdYehJ0cbSAEoqAcfx7aNPndjhUKtMAmhF/OgT/FfXmO2At4vAlbzAdMjgqENMQj
in1nfOsUd0QuYto/ccSgRbrk6iE6kd1qkcWNrKlnznKzjZ7+TWcIZwNG/oEwI5KbVRbhheKYgKtf
st7YraU3VUhbdEOh0vStzc/snDf2V5S09FQ3GrFaX+8w7IsfhyCAR9TQjYBnygD1iJVttccnQ1Nm
iQTElzn2TOl6LhgQXb9ietExoeTKiNWhboq7DPyxwPvWPojGSrFmWICE1yGumdPiSxsFnsU7tQkc
Xp3EY+nDa3DBVeFPhCbbyJZxqJZbYH2x1grYYZu/F/vAaAaxyQY2lKS2fbn3w6pwo/lOVzjnEDtU
gF9y1/tD/bzg+KkUj1SJMU4W1IlxYD9S0M4bYlB3WInXEIn/JOxZuQbOnQ6ibKoFrtCGgF2tJ2VO
7e59NgQUMoHEMb/7P1W9gXggRrC55spAJaZWRt0v3zlXGX6AmRTRKctplt62WMmqSATwtI8BlTBl
ewDr2M+XC37F0UaEq99tk1F30NWk2qY5t4CL9PL6FQqGFOIrXelqHjH1KKR5jkE/92T1dMqRoRKT
YUnYb1+Wdlyt6YC8ILhoqMbqVBnLrOioGReAgsXjJvmNty0iI+k0N3fcGwUCDGk9jo11etMEoSam
jfLEzgzQ+NUJguwAFm3MiqDhZdslIrzB+Fg4YCFJApQ73v9fDMwvZc6+e0TgQe259oe0QsHL2EkU
93TUiZ0yvmx3SH7tqNMFksmM17JtI4ZWTiWurzOheNNUI0UciiNmB2MiCUV3scsDINl9uFCxYFiD
yWC2aiIHfN4JPY31wpeR3mLkdrObHFw4MvdnQs0SsL4g6lgsbtg/fJZtNAVYNkc4XGhyMncRGZCV
Hs4BsW/xC5GAzdFnI4Lz4JgYL2LGrGtJaeCotXL0z9GQKJ/KiOcbRU4mi5FKdv6xqz/Gqiw793yH
26bcBjRy/k7VqibC2xy7/OKD9r0wPIxE60UULZ02EKnhgvu/kEVjsLNcgG+O0sVWIHaRshuPu5s3
wu4ip1Rn8xsYW/jy096Bbf0F4Z2Qthwb1MRXjfA8Fa4M6MpJMUXzNNljzwG8suzteaij7kDalbOv
BEy49fwWSqPT0mJDm4du5FExKfXNQE6wkt5JWM0navMs3dsMgNGp6P54uyK167DkD8bqbVFGuc6K
RnC9HpN/In4KOcYVryKhwE51t22yWhfjklPjTRAGJXdtRClK0QR46222bpMkkUCECM/d9tTlC325
JHT1yYg2VGYsLKHsMcGq7Vlu3EHferERCfCoH6LmLjfCx6G5uNP4c34APZKmtIIKFSQQB/FlO9g+
8J8MA7FfL6Ilw3+Jg77Wb6h90TzRUTypAamd3ToHjVbOJ0sKovBslBEAw4icd6xN8YswGpLdRXQE
YmWvG7EA5RvF9kpvmAsrx6lWCFida9S3mmJu6um6vzEE6GyEmoW87kXrjAFoEti57lgatUzGQJhF
GWEsFfjuiTawrzfa0u54yL77hDVyKu9O7Q5n1o6ZEUu2J4pe8Ww8ksbfZgzWQMaqIFvOIgHXDpyb
HN9J9vstlNYGyaq8jR9EAR2pJmXUkOuwNCTUqWj0VL5D7Ena0WD6TUD7WghWY4nJsYjWNWrIxg39
JhRBzCgzOoVlT0Hf+STv0/D8lokqXbm4UEWyRVomUerYSLbDej8/eU2+Hgp2O/BMXXljKOc4G4Uh
y8o4A2cxccd2xY1j78Li6hN9Us7+nxY87VQJwZyVm6OR0QFbTcbycq2L7yGsrlZsnyo3cNSQGmZE
aJ4JIwyBNmsCaoYPYPhnkgoQnPtOTkBNpxOg2zy5oi0nKrurQGb/ClrWPZHMAUorx2vJwY+2HQV0
fBIsKQRLQGL90qfFF7yHBQBGehetDztY0UYB3rl2Pc2EqHYofEO/AKjj0LPDQUICHtdw5MOLqGrr
2aDzRXCP2ZNEQtAxwuqQdIReZHNzP49d31DsLn271vys5PiAA9h35HiFeHrF5PfHTDeVO4yzYapb
4ehoCUtVCANygQ+5P+TEnxcwnEod33dz2zhZgyBfxAbS2NONI+2uWcrF0Y3XWJQZh9XMtv6+KxeN
uY9KJ750iLYS+nwdMsfK5QE3QGAtE1Gc045GKahkMlE2a66PaklDih3c+DD4eht30M3/0nXMMg+n
4oyM2MJtS/pi3Vp7c+mp0V3LgMpdPaLyfspFYtahbk/mnmLTWgWRYj+kjMvPST1qCesVHBehcMdh
iMcJznBbMxoVOEOM76X3OdxQqSkGNxVsJN87nMbLjUG03jAXQff4fT6rCNm39v3XBy/iMES305vq
IXlQAY3jcN0tZfph7c11ltRCPLIesckI0K5Eux7eeS/1leW3vCao2ZukWZQBeDw9qF+nBVQfNhE1
sisXmEDbwB94FyVmFwiwxcWBUVpaUJXRMDXzLb0d8vgic/JYBsOsvg9l1kCrAUA5YlZ432meZgur
pN8Ou2hTCriiXJD0Z7oCmqFRIUikhMJUp/Zf6NI2im7MZspCvaljWOKo98Tw5E5KwHTXlRUUWJ4p
9jRP645PydN3aP6m3QBabElQuRl2KXVqvArSkQqaTdPaCM96DEG7ziGqtThmRV66+R+faxZBvYmQ
bLVH4jgt78c2vkBi/AuzU2zu8nckPxKUWpx/s7coFs0Bi9JAXtYuE7cA2ksMD54bMYkN3xYoYDn0
azWaHQCcrR+oWJBlS7coxV5sPRph6glaY86n+YQ0eakC7cR99FP2uOgQN3KNhXwKzE6/SoK8qAj8
FuLTLaEe5XDXZPryNJUT4ahp2uLlOECSEc9211O23cFQMHc9TOb9RStpS/E0YW3enW8wOtNTfIRi
p220EQQPdtmwpKy5P2LVYeNnTa0kGm3ym6pkiRBCspDVyFkMKgkWDa74ziUcm2H0GMumWwJw2QJW
vQaj34QTusvfswvbloP7XMZlO808JXz5XAUa1MKBaArOTWXpWb6UB0JMPX4Z7wRA6E1IWzYMDAa5
cuNFsE9VGdE1bK6hAx9unmEHhd4PaCRoic3c0GhBcz3fWb2cjeqG57EEtokMVwKoXhdBYL6NfFJ3
/C5jlOqzy+m9ASqXMr4rLvXwVrSjvyYRcdBIpYLmHQn24ushvEbPdXdNLipj4xVGySFKdxzFBqRf
2YS8cDpgg8MjpJ0/LSP0YV2n/puMy1R+1jHppYu+y2P8TkeieoPcCkDE4BVQjEJbc9BT09FB8ZzG
tQLnWLHu0iPydCO3VFdcQBMJNIyGK41/WJ6Dny4Obhx2VcjEO2fksriV6wm9R8HtFU23oiqTEwfD
TzOegbl2OaC140MiowBYIUKH0uT3Iwdg9Sr5H6i8YhJ4GqyeHwHlliiTA/a4aQjDUE90ALVoijuo
Cd44z6mS2Fpc3iNxfYX/n0CFyuSDuAdmzsnQmzd7ANI+5Sv46wx69NG2MdT9zZi6wUKlULLt+q68
1u3PZGB/YMnvugEgz22YNOXK/iDH2MG8Azb5kPkGwtVrQ118Baax6AmsoXPw0m6/JNe6nB6Z9rdO
mGNPewL6UleV0j3+Mc3watfFqY7vYbQToXKajY/vqirKQlSACd68F1Mvv68Hr7D7vZix0zKgW1Ea
D1aPhWtIsAMD1sdERrt1+Pkog20A4IET4Sp5aXDyn0e8PdD/jmg1pP7+qylCpJZeAATZ/1YQF7PQ
+4OGtRa4aEQ9nJCujVR+qzOzDdMt2tUAu67m61/WGJ4vf2M5K8Of5hPfgNHV0HYs+cmens1sdmar
nHGH6iImVP4S4+rvb4oWyT2o12SuwOAyWV9F1MuHqouAUWWdSJeYSPBQnKkMaSqP+4G9v5N29Du4
OQ9Z65O3RMid6l4+hYjjDPpTaGEvm2HUqSDz0Gdp5JnKfRGJyVbjQpbLjceHwXDv6RjKU8u7fRJP
oF+/ZLSs6sn5bd3kksri1jXKYyFIl7ubW+I4OUv2IVFz5cXCae0O2JPoqP3crxx7fpueoxr+oG6V
uAWo/2hysKZv8eF/tOVGyq4lL49RajmHNVv0N3+nzA5CkC6iy6YByPQnx2rCY9F0YE3w1c8ii6yV
k/5IZ3hn1Wbf14voeykP3MbR5pE7y538gjrtgTsfAV8lAbh7EhPKaQCMoTs3eBULKWwmOr4rIop/
Cp0q6NFLFlT69lVx4z8O/abTRxqp3tEejurbfXWjnebex9m50ihZRyn0+0rOZ4M42dYFybFtrQHZ
EohOd7yv/HFENsm/u0Y06Xm8y0oX0E8gX29BGP/NT3XB72W75N/+CjlTH2Zm/0wHgVI0dp7Eu2yi
tXWuGbJJNXndqe4V0r9363OuTPZJfhOMxvV0fBhdohTC5O+SBwddYqF20G0A5uy4J9tzYvp92vkC
0dYX+ADywcdOBGwrDCfgp2/1Do6kuzVWE+D4+iP7uUDyZMgg6CL82OYr+8InTqpuCx6e4Q9LgmzD
pMCcGHEuiXDYX+FDQZqmAOJQn36Dp+p3KX/TpKfdbZEyswcQQEhiRNfzVcWtu+Gu9xrnT+hwxuu6
F9sT0YOyx29RntMil1D+NVirVKwm1HmzY/XGnLrG6dm0xGBbuFe26pQ/FgF2xMEexETswcZEsbC6
7gFln8Y2CElaG5XII/JJS/dNvZXBghaRioNw0Fg+7/svLh4whyc3i4pusiUW1ag67pzRDqCq2teH
vwbwr2bfzPKllmmWg3BmEJ6bNY9i6WbIvDlCRU5srzEy1WoeAYVYIQUBKruBCwXi/wCmHX07I4pL
5olHVUFDjKDZRvingvNy+ZdbDLw5Jx8lkUVEmlo+4UnCd0zeG+Rh132gwe1RDEggtHf4lYrrDGyS
b8nLi3gAYMzCoXjGrKTbLRVGZ3ld4JxmyyOYt9r4z/57Gde7kcqWDQxfpUdoB/VMzOfTDRcnTmS1
rohc/IY9M7ycSqlZoNujOCdjd+eLPcMD0sXxU1eTWIXf9acio0jkGNN7dkmZd25mnLSERH8xES1I
GDHxD0ImOd+Tb6mO5lNVXR4LSAkrgdy/Yug+pn4/DPfDKb7U5trfo3wmdoAxDOTupBUYl0PsZeOU
g3phny7gMJCPCK7QpoJlqOpQDIJOzuJGdKcXqK66P0H3OR8n8Gb+6/+x99ea2gg+Ukoe0tjbYovP
B5QddJxwspOG8HtktxQlGFelMY7CytnozIUpj9otcvKNBbIv+qNkdSQIy0UGJ0xb/+YsBZS4kzH6
PzS6eJxN5CqRRlXOakR5fydwd9oR1BW1M7gECJiIZhGiKVIMmn+O44bHF7qL14bW5tTM7x97YOld
+ykUPJxH3STkodfJ8l8KrJp1EPu3p9gUe1hp5fVBA4JpnnT+eyUtWVp1+EEnBAaAS61j/EKg1EUp
sK0tVdXhCvargb5wsoav42zXPqdGdY/8sJv1l66bS2xwpCUh1ECO0DDsYhUgSHzKsvCiQHnyOG5/
oxdAo6pgsMb13ArQNV0LkZxJE0fGP8jRx0ObGRwmZQyGXCIx4Peu6/2SoTpIbw2AAY5OMfvKbDwM
/p8vVFurX5FZHTmYRsiDOL57Cr2XbL6ed63V7TcRmORztW/yHLUZmlH0RY2DZeKCpS0lXz0us/TX
p0oj/c9stdM4X7YqlMU6LMRUAFOJfry6tzwJxWmRG4QqiG1RKgGWIFMOR7C+B+Veb83lAauyHIdZ
1PXfvcFUiTxWjZUQPcxdD+rp9t3ekrsNiW3YLRIUtnBmK/ariI3XxbGHTZ7c09CV+OXIjzqEk++0
I554zv50nRvU511CbHNuFLRbL/SIV611lL91xiH+O+YNDLxoDuz43YAv+lX853Q3VhG1JbzLnX+l
CI9wIfHmTcAVA8MsfdFDQuPV0UHdy6e38r337AwvzcFXx6OPqAbI4+LYPUCEhwjLC1fJ9gnBFWNa
Kif/d0SnRmZXDU62Hx22h3XHmVeIOjRc4PAmXM7oLw/cj85rW9MWwHuWMMydid5Sf3dtUeJrU9Zk
PMqj1nz0WPLnbc5plsxbwP+/GwT4DkuE+ikAu99L2hrG9RZLpvLFsId9LrLIXBEe0SKM3BOAWgtG
BpEj4QCtFcimxcQHkUEv6gYzXFphlPMu63h9i9HJ3UxHxtqQ6JhdM/PI7hkWWzR4KNbhEM3bXreS
Rc4JjevPDc8InI9V+6UYwxuFz2ivSEowv88iovZ4OOqNB/vbJJISVB1In5EiyWIrlVJXlLRWrFwn
ZxikWu6U7JzNiyGnIN2x/idGj2W2FuR+ADgXjDTj4uNd2E3PDk8WQBbskkt9FPUMdldXKBzkStfz
YQqqwamk27IJ5tMyzTNg72gQpUHda753RmZW67rz4uTCU2y5tHutN4vDx4FCb70fNEv6leWh1Khl
MnCkuvI9FjM5tOlccwspVU6diR2vXRB9pbOsM9fh3++ext/14gb/EmTiODQzSsz5qjLIgP6yuJlk
Y+NAjCFtynbbwGpUB6pgxwBB6gli9FTKyjQbGdYnssNnJecd90W22K5YSntanlwDuBJuxI2fMbMN
kBa5bg59br33UB3anlWYnEgP/aq5XnLOZj7E+JN+M8z3nxP7oYNKucx5w4MPHnrPrkvh61cjVOnY
ZF62rgpfZAaXCmcPY8B3rzDCF3A75o0TJANo6x1XnB/+6eJGfwouUPZifHXAv0jvbEVhjamJ2u14
ROY9iXaQKCuLo8R7f1NxH5JrSg0Y2WRvs8D38AhcQQECPd34zzVJMh/Z2shWBChRXhPGieHuXNWN
Lhsg5KM7yYvXokcGkUwec0RPpL+MNMAvwNQ7naXvMqrhou7H/YojXTIYvLuLQjRlhna5/6wcXH4C
EYt9vHk8RPLwazQtKTVWF71W3otWD7YfLMUS+dcK/yxadhdFUt71X1f9Fc8PpCVAopk5UqGh5oCn
xwZZsNMdqIWOriQ7Jq92JQyg65qkx0Ljten4eNg2FGnwTWz2wxz5GU3f3cGpitaTE7MFwhjQQG2o
RKAkCUnpMV4QF8qxWUni0tFqCAw/tQJpXdDO4iKjendgDf5aqFqvL6jM9bRaqi5fj9z9TtK+UtOe
wpJfhER5kTZqVwK8sY9L8ujIqPSyXM2TO7oSh40NIIcPUHYNToL3yNxZBhbMZmW+Vou2GeFWzEsQ
50x3ur/Rtkqu4E7E3IZmDyOqvBUggQoGf7+SXR+3QCYKcejFzcLb/YZc1kZEFoetSzG/mY0Q+tDZ
mPecQcJOwqNh6hUq2RTmxz8M777hVAlLJJwqxwPWNssp+WVdhPyJ4OBDYS/J9sjJmbaj5XVzRypx
lrQqb0KQLNULHgwEB5PSMB8GWoBgD8SXPImnxbsiSzZ+JXHIcnvetN13Imy/ZkzUs83FbsUpc4OQ
7DLOW1SjRqKrRAI3fmXraTFLO//2D8oLho8Tk1QOg/k4nwaJMSbzfii6Oe4HqwQLYQaAsxDS0RIr
ACxl2Q2xEhBHVp6ZjuSJ7nUsXQiUVPMftZbDOzljFdUFtftYe+6UyoR9kngIVq9zaQ931WqY2c1O
+hOO09yPKifcJkYiDmUhzfmrrdYuheegl7v/L+cZpOvyeFZu8eJf++xOkZGDWqODa1NLwIsQL0+F
AyiXCCkhqjHaPgGAlFMAkz9WuLDW/0NYAy8CSdez/11lO+qHapreuIEv9y723zk6LdoflwPxGYXk
0iBrlD+/wFtp8MiLwnL2eMn9POmBAULQ5CJX6sIQnerX2MKNmJhopzKIbhRhC7FVbHvdcbHSIZFN
z8Yr91ovZJzamfj2iDaxmRZjU/Hp84MYcYWUA0UYnJqr5oXhZ+vH3lHjh7efawhfSfzxPdNZliNm
iDvRunRQseMx1id9P5cpiHMcS30zWBydo8IIhF3JjC3VrwlXeiTqNSU0uxju+G9Y8w2aAzdBlgp/
923559vYFGfRs471aBr92PRErPqqnPVu5XEnLvxTDMcg/+KPmYH7RAaYRjfVC4uIMp3k3fyGICQI
nbK8F5U/oGAGUw2TEINABSWbFv7fiPz3J7nOOEwCJ1vv397Rwhf1h7XVy39N7PE5t4ovMt8+kgf8
003SN//4UEzkRrDTwriTvQsbZNOHtAzjs6eVRJFFwPnwCqpKomnNVQ9Zc7XtVgwxuHAYWJy9Q5RV
Ds5CMNNIcwv9RDqBvEYywhdqIo0tOcxuLsUXVHT9YZtGNKjBpoAhnyFnjnCGc4TltC4QGv0UR000
nJmjho0J/8OizbSqvwN6LmkvlJobgXLIV/d5bxQa+HlG/xw8fqkwjsEzTEroHuzOlj7Dkfbx3Cqv
qhs5TdC3hQdPF4zpCVx6PzY2lHdb3Vhnu+Q8TDJJjNfDJlY/0OoI804c7nHDYbIz/jnmGjINwFfG
0caFfnVPG1F4Ql4bA76ILJOrMXX9QYinWZs9KbOq224d3FcPwiaGW4f25P+CBvxkVlLQbu2mSrJ8
YO8DkVK0Mh6ZutmhE4s/fMzCCRZqAgPui26Ai76Sea7JtvpWF9SkQOugH7lG4modkmCb/c0rSjth
B1b9H/gB/Hh5pcbTvbFKlqL8yeqKTnPsZ/wL0OU9nGHfSiItcSAykwC1AqXYguV1icwWQk8aPzVj
zHSqTdO/OhPbVcmbBvRLoC2sIRlYA+nfRkq8d60/VX3vV7Ka5xL1TcPNJC7vxslqdnwFb+wrLiWQ
Ih+9iu5p/0KZuk2seXBVJ5bMeB0dpI/V0h6AEh6KHACQEVhamFE7CRnbiRgY60nQr1srmqSnfHn+
xIvKAewmgouUA5mgk8ZFBcODv8SOlJTCgFO47mrAvE/bMF8ZthuHCwiYbRv+y8IjdJyMJsp6SM3T
WT5E0yw02Xgz0edbA4djnsks9JwbnEywmrfeivBtYrxG4NrY2eOv45e5Xt84Jwcx14JWAiZNtNYJ
PU2LFKPJm8qyyC68g9OIR85/qRjlgOnP1D+y4sXQ1SRPUQnN5Y6KsgN04wc7xExVrFKEVSlfmRNQ
JOg4bI1l/fF7qGtrFeJpgp9nbuqpW1pND0noY4nOJIGXjLYJCjmb5cmmCBdHy0dM00hFhB/WRxSc
ZW7oT37BJ4FXMlC4ihKmxy0T6xEY0xvBJ0Q910PbhwcsmiuXewH7bzH4pA8YjVCrMPTl2sAsoky1
LFCHdwM+yfWJhNdqRTXHMSGV7xQROSr9v8P2XAL7QzPNMOb/fjOnw04j7zLQx23eU7RCjZ+W7b46
HM6r/NGcEhAre8zVlIBzw11ysOxNkQCL5H+/q1GkHx1NKbWiZV7XkLczwxD7HTBt7R4vza+ufWpm
5eHXzCEYLYjWGKsULdHFEtiYEM8mqwYODtpLjY7YP4FKn9utnuBazad7reuSaLgAWvMh7CZ2OAOK
Hu/sFkZ5wywjMzaco8lgNRvlVO0Ls2G3k8Al23uvHco1BEahzrqz+DLkiOXleSdLR1FGApUMJgjV
FI/ahxzfHjLIa0oDm+yddCdDfVuX4Tosxex/cgVa/wo76XqKQql4OFjhwH4CVlcb5+FdGPlzt1Tq
CEuQgvryEDpBQbLF9AasW28XxoJ4j1PU74RpE3ouGIuoNAivMXTzc1JuGrzoor+4nFHKGJM4M2Fq
Bh7QWXIkF/oBQO6U8IiAEXKtX/rrIKu19jqbfWcp/C1MgSMQOm+uzdos7weesHXjFRvJPmvFTjEy
qcbDGN7RyOGtOIGzW6S2rXRxjmVNtKy8NL132Iuugo1fz55/oaEwAZjuxvcqCc4Nu8K5nd1Pi9W8
6Gujd4xiUUqnPvDs0FxHw2ZGYMUxpzLAqk1l3Z0JoWEk7Z241EH4sXdwJyyKrZKCZwghvn6e0bte
i6UV620Ai7/9wTWCelTP/upRhiw7ZRvs5bSmAH38cXLCqckuDfg7rw6zoI0NMCaPdALu49UnWFsN
Krue/dfLxXRt2LQUiD4kc8HMJT3fkzONo1hU+U3WvqezI9fQFhBlSZDmdFVTYH3IfmwCnggoYb92
YHVt2cqbiHav3YUh/9zPRqy43XuJAAorozNwQBe5M0bKaHPUTyFuln84cD68blMuF5MDpxxK+Vfi
lh6Ve74ffTz5vNmOaMBy08R9oXTDIpt5m3uKmSQDVylP/tlXxdQ5JlyU+bM/I2ZEuw51b5+HtLI6
uYk6Ghupop+Q4SuD1e6O6v2uMNWkoitxJzfea2v2Mjmxb0xEiOrwo+/xZaEgFFujIBhbbSKYaArT
htdZpMHSL948g5okytICaz8O9LPgsGSnp1bME0CGSaerVaMk8/OAJKMcqn6iVgttRpjoLd9YC3zP
/HyIX7497l839jRruydccCoVnI5VsSUBF4vT/pm6ZoUfAQGDRu8sFye060Pgo+WnJyl6XvK4+1+E
cqexsuAOgi6/s1eI3YWzyOeHKgSULpkNaA1cjCDa1bF+rkHkP12/18iW2AiiPLEHLAmEYFM01tiE
uP5bmloLxMF1hnVxm6UhRJDUyWbIpHFzTym6ZUaJeI7u7K2y/1jAv90cy7zhqjNq2ZAuETtq24EH
Bqc8z6mbjz+RXZ79nVhZzDY7rh6mvCjFDuG8faYSIFyGyUAVaTQLpUHfKeXfmFSPzLIODcjhCDTy
LJ8KTFQOhzQ35o6IGHzZa2eVd3oUOHFXq0E7gZXI6kF6EQ7u4jwNZ5D937BxQnJVDs5rff4RIgze
1jwYF6F6z10gicPXdcYZEdcEgIrTzm9bT3XZOgL/pryTFhnqfVp7EMV+Cb/p8cOK6AoACEFpc5Ee
DsgKktItUv/E9o1Iu/dtt403Qm0eO99t+urvqfMpM6HCoqPLkotegNPM4ER5dyBV+pCnRQgCg2q4
NCOCDudHv28a+go26jn/xP6alSOhXNr43b04vKsmbrkC5MRG08QfhTYwKNkQAmimBPzSbR2ZO8MQ
2Z13kXbnK993x/xZxdnmms8Ock+FUyXUTlkDYNqtkddDwNsuG1Ej/v9zYmQHANsEi6a/ukTRNZn4
2+zC1iKY4Y9xxThmhsLRle7EBGLTB7GUlpAi55AjtmXQZSLJKHYelF3Q8BO6mbX5Ucwm5wpKdIMD
L4Wmg5b1vDRxwjg5h8aM2NfllFdnGFM3niSY0/v/EqK2wTifcz8aFgCdwJeiIV/gEwT/blDGUzSQ
YE0F6MTRvTEq3oqEV8vzi2zBqVZ6mb22qJ/eZZvzSL95z3mMJcEDBVuDKrZuQQjTTXrg1yZJCBp6
f5SEKVg+Ofi9KOWmkFvUxfkZ9UEv0JJxjJlEk67WXeE7K1TC8eZJtuxg3sjDd28t1yS4XQg4zqOG
0jP0DZgbTtljXe0B+fd5ZrBSdHa09jHITa77iWI09pZDQeTOL+gqbyFdSr3BN3MCow8V9NXYPyMN
9o4vw1ZnPt6XtTIWRIdz0B/sSGPKWLJx2YtdQwhoNAO0HwqACbxmJpokYmRkKB6URzGmCcTD/eVG
03dXtJ1sNfxFkYdz5iVdhyRxXfIpR2+fMzku0Dz+JMb5goAUvj4f2oDjkncbtnkFVWG6JSMSf1zS
JyW5wwO0CZn271q8zMVUPIuz+PIod7KAGAsCxdj6LISWbgGT82AqxZ0ynthFeRAe7nRXaYvRIsE+
e/cuzaulp+ndY8bUg3blxPZ7S9gWUjl3Zm9fkCmf1uEQg1oTgro7tBMIEIZIa6iT/zras1t8hDX4
iors0ZTa/YNNm+R3XO7hdBetTax5IS21P4v+njSaOCRBTvNsoMVtzt0Hm97N6cFJzqQ7qVT/4Q8K
8af+APoYeWgo5/wDCXIx+2zYspYsY2r27cah33ZqbmJDq8lWgM2HYG/lhHPzwgA6vSRfXZFpuXeB
YXgmk+lR7F6moyGcYMZSDpBQhD69x5T9qH3R0DiIroMMPAD62/tvMZQNqZ2agZyrGBKZDHRR4CtR
jTFAwHF5Z+mb76OrCQhGydbXJS4fxrWpRsGanL9KMk5z4j9bsDo07Ft3P06rTau5mx9YYZV94fg+
k/63VkGZN16pg0rdfX3f9kxDGQ4glunteXUp9HejsBbLkQ/f/57PnkAfJCauI63vXQWp6FDslSbY
SCogcc8PnluCQSuBgxcjQgmKthUkD+6/MOa9Kdnc4dXj3Bjg9nFGbtx2ultE6MQ8+Wa8nYAaljap
PSELfS2ftNMXNxrELKrKleJgNw/5Dtnd0+KmqVkcZwMn5fEfRZXqer+A4EW00IJJoAf8MVr3Kmaj
OOVY3Dyicy4Kvye4dbUf2EdesMj9d8+HDWLytmkbCZqWc4NGmb1/hsg/WxMH0l4I8vB3XP8Mw7Ya
d4lxz0afR51JAIno31zmyyPAr0RSlgTl9qiLgJFvg0kt/HUFvb0niwn9qjrolQsr5mLGtIof4kOa
/bPGAqGb2+oOQ+VzLvDGKjkyrFPfyS925ohVMv8DQ7QBWKJWB2dV6ULyvsLL+9xxVqk6to/RqLbK
i2qv3Xovr4DYXG2YllCdobKREYgXwFQY00mfU18FysF9OtRUmgxEerW2y6rNK5ZyDeGN2w4/u2wk
1gI/tfTVnWigWNkp+KQLkrQZ4CfhCwKkKlS65vl9qetGVtJMg3dwuFYHS27H9XrSToI2JXZlgxo/
3+rL040y4Zw/7lpZldnlaqw66Vx0h1TKcKAQdAjOdHPK1l5EyLXqU7V9o+GRPB6mVJULd/WgHmDt
aTO6XtEKwKWzJWhBWigLWs6dnABiWaqqKGHqDjIxUrWh4KsPJD28ChR37refDZPipMqvg/UV7Qld
P/IOo2Dg44KWOOLn32ihrZ66CS6vV9lGIa0oN/+oP32GU7+F2pCyWhpDv6WwPGkpOAhzwsOaEHA3
/um/sD+YA13UiItvvsO5VVL42IOapczOk4uJkq2zh7fiGRu35cPuLABp88Vk27m6Qq4kI0+49IDo
ikx+Ri10leztXLTYOP54G6r9sSKj5/ghIDw0AbT4da/1wVxBKbqbZG6EZJBFY/XLLwyIfr6siZVt
rZ9nRWpMmsNGTtGNAYB8U/TCjxlN5OpQLLjAJ24ZCCkQmwUOLdcce/d/Bnawbollmhm6kNLqzv5c
25kxvmfu3vlhlj9iix+mDjJ+1OsWoNcpVrKYyv0nUNlEW7L7HFNeF8S1C42GdabO8xhuELWmwz6u
n5ar4q8bEL/uEHhcOd3z1o55znhNJrhr0G3vpAAC0cI+wEhofMQs0nv+3sj07Knb9IjYFhiRz6up
CksaNVbvHL+kvKFYCOdaahWmncpKbcod898TCa5SayYg69qsNShkJ0hkH5zs8AErQ5gbqoWzm7Q0
6zs3KnLkpLpGzCfsN+u7JFK1LtBoKDwm/knC2bq0DNYaPFmBQLqt57UXGncBowt4uFf259Htkk8R
IOQ/NV/kjetVYKLxI/FULVxtG9Lfk6K5IY9BQw9gmya2d50knIdRS4vHJ1eGIVTxg/shLYCIrm6u
l5Vjz6PxFiv8IkU/csbF5XJBXk0eOobcBfhX7/xDT4P00cZYalldj6Yv195qsLm3Y4Vy4oG6mH4Y
8JbwtnqYdq8cXaj02zkumadrJIIP9HpqRQfGapRgBNH783e4Uky8yAHWyFezs9xvVQy7IGxYBpJ7
DY2LugavUtfkw/waQh4mK4H2I/0yvnitP7fLtlLUYYyv880impPBK6mNVkiZdJ/T5a5waYGTYB3f
1XejqvJTODQaVQXSHEDeHB+aSXoX92CYYIOCUlyc99KByav5en6qI3M1Gdz2477A0v99iIu2KvSD
3hC1hu0ophu9F0rgCfD1d5Zq/ot6ghcuxCvXMGTZHIPpMhQum/WeJuFdth6kX20ObEE0Czsjjmh+
I1/dCVimYMffiA0qKA8pSTbULmr4Wq+Ii/m1xQcb3lKB6H8Z9NFeHN4sdS+gzFC7LWBF3hXaxLix
fazPBQkJ1CpF7zR/ZTgU1W14FnAsuM8WygeylnjMowr86bOlCScIN/5ZYokL4/JfDcnvkwcwuknY
wICQEaNNmJKdc9vfVYy8S4WvoOUEFZxjNlo1/JLHz1y7Ed67ksDH3/cWKr+oIr8cwCGkjQQXSzW+
vpxbn4kVpx1WOkmo+V1aFhuzJeGigXPwqg40SHCJjzezjPRRQ7kneaRBNJSQ5sgWA5CdSt8W3uFJ
YrKGeS2YMW5G6mAwPB4WYRUf9qC+3wlHzptlYw9M4BTF6mmwqzutRZFyCWCdrR7eta+VtzmL3fPf
+Nk00kTmJ0lfa/pyMzIAbIWvTGf+AvA1BR8L8ufzDak+uvO/sgHLLncU82Fe80Q/ZCFlckI1fedN
Hp80MlAXeItUxdEv1VqzEtilkf6rZWWhn7hdcAIskDOKe1BQgb8uRWkWbEJkpQi0rPJfeGYAuyBA
1s3h5OMLtJzDyv3VfLpj3wx6lj5ZLSKEdS98pnU98ELORQ/FuedEdpSkkDK3vZuZg9Kt2W5Q4NS/
LkQlCGiQaMZd6rd4sD9D7UjsnIO1IJoKwHoeyE3CTwyrNTXuGrsdR3XT3EPBurhsrSVlF4aWCVDZ
qFuFzuqWogCrlOe3oI8CAqiPB6a3qRsmQKwTaAttJFKccdalM0FgS2oevwEvPMB5Er7at2aHqF/u
akA1+lW6YvzChPhrrScC1T8xl02/203Ikcyp7qEIXQqo3xuPVELXdjlozPcMYA6AppRb2TWFdBKw
OTyz6orHqDsmhUmzMCdtOF/bR0QPJzkNnx/bTgXHIjFiq/nocgv+GM0Pu8haaziejusT0o0FxvLK
iJ3IOFlG7P5t9FGGKdde0Z1YelBOCa+yzsZ+9nD0hOIoES7dL3nxBb2By/1Wqhm+0TZptvNH4vWo
xmTrTwAKRY8pUfFRWSMImeZfDuHTFvFlp1wpNeNtgatIPnZ8uRP/r8TJFAi/KGauhFxjCmgFLCx2
ohNvLOGvOLiz1TEQGWEZNnIGyTRXUmOHw8OMDlUn5v/x/1itMTT7YC2nGYaHQasDV1ZBeGTAcERs
yWfYVcA9UuJaBuHx/k/eph0+FTh4Vv7a3F+FljvwAc3IBB6JNWIP4O2AGPW+qI01APC/5qqXy1Zo
caxW5EfQmW4pA3ACU8kuK65oHMJvtb56r2mwKS2h2LUNgyOldCa/n96Z4nKLqAxoobD1gUuJKdWB
cBGFlDitQ8WWXAFH8VYvZxGfovix+IkIYjSyAK8TDyfMGkIN0vy29NxU/CQdtQo5XSyTAEp5zzwj
JNpPEt5Tv/q+X3OLyqmVYE0ZxPIhjCOM+TOgiAKdXt39uCjp3qfekQiDwwwernIa3cdbOeVSwU2n
/M7eSRvLiUpt+DEzZz3mWdNysyaD9eMB2dxbRpA4v77MZgdLcTvBRpR4Mm8XKWo5DYBmSTvIyQDW
EKyqMNN9lGIKeTTpvZo4Ax90FLUnYuit84k61gnVDX9QO5cEjijj170octvv6YAo0HoCEj4ARl+b
r2Q61FftgQIT7/ZpIf72sxPLcr8dR5tY03fu0cNUGCd1q9KuPFRoIS5Sn6Frrbb66OSFRcKPSvTW
+QypubvdcQddQGFZoW1E99zYDRVmalOMIKPCVkrit/UiSnXEvCQefKyKtvtiju8ynpnSH4UJmMiM
2lCh7QIjjm0jMqoBW+aLQHi3c+kLEXayzFjT4gDRW2KC7P8j/0WQS+sLSCT0UlgTW2UBJ3BZhlra
EhnW4AEthkXepvO3ed93UTLVxrzggpvPt1kmLi3dj5W6UXRAU3P6HgXpqfwe7dKT3QKPr4VZcGWC
aYnUTpZ2c0mapsu20pfUvgW67F3UllX7LHOevZTN23G5SwluKwEfyuwl6o9eC9/NYXKKjvMoo/vI
EW5Tk72UjNl3yoj283LbHiVMy6YiE2ksJZWWCFbDC1z7kpAgXY47earcPbeoHnrSUBb1L9B4FkqY
xWDAy/EG6iDK3o37iQVjNIzd1oaJcyLw1kBc63eKlXnFZZLxIDc1voHX1A/7SmY/oDaJluabyviC
maz/EOPc/9h4TQb/WmWim/ugZHNSvlzBO6Ot82V8g8uOUR1xNteAzUSMrehGlM5iBxCRl7Gu3gGk
DLN3nDgUJIbJZr1CbnEEHn0RpsJqiAPqqP8yUZKixAUB0NZf1t+6NkkjoXqQLHx6v4gYby5qc7e3
jLHFh+VyweThCYV/F1rw+LHuk08nkTP5pM7408eLGLKHPskTzaeo7JTThcYakF9/zW+/qv+lTy26
eOrvP0C9sdI2knaGYL3W1txzXj+5kc/ma/s3rrjknherzLwToQXLwjYQTTJK3i+fn5xaQOdCGFNI
MGAXVpKRl8fdRLSQVg3WOTB8wG+gpERcma+YoHPM70HwR3I7atB0KfXh7aFmFYZJC1bzocetZ59R
ueUL4JejiAIaSri2ND5bPV1iklJlP9cKZghn/C3U3/RPgsbUHl/PISyVUYmL8BY+vbol1cL1v713
rWbHCSLls39lpU5VAFBpTxrvHi1eXt7SaOdwWBlaPDqF07rZxJXBucdz10sLWYIRoaG0Ow3ZO+ha
BpH3FFyajsc3EByP4UdNPOlbTuk5G8jFua1+0jhT9+n88b6chrEEhO9W+sWOPKk95O9UKoXHpOQ6
xVL80s6K5b+RKSplUeYCfDq/Afqqv12F5cRzEJClmI/ohvErEDxe+kxlkM4hMGl8ZP83IPYmEkC6
+3xYrEc/CdPeiygNCDa9APlEDo54ShmJVGC4y9dtb+lrjffM66TOdzh74uZXPpMPUCt+z7x2sFiO
rA4UJG+wJ5+JjN8zww3zc05haKwls4LANQd1x2G8xBscsbohOFD6u6w9AFerjrrsxaZu5OVHqEAa
rLs7wlHr0d9lc7qZsfLxg41rY4uzNlDdLXgpqz/YdHxJ+DQjrJNs17mqiFjQQ268QMky5w7YW4ms
x+0KSVKBGFtweR76HcLUBKwl7pLgU8P+LTCsRyYv7jqfZAbZfjPgTn3uKB0nZ3TNzbS3rM0UPp0Q
4jpMNgABQ8sMoDZbmnW8RmkLR7cyOdxBtlaeMxX7J8s/N1Fb5qxv/YPmY+4Qga62WYEEWyV4L3WY
SqmqWH33+cU+vN5rhqDs1aT73UhYC7uu7thyhWw7+br+bwtaCD2QB6D5TGPu2Wuq5roeGDci+yca
KQ/fmtMtCjDaTvoFmqAO+4WVQguc88wKJPRdTvBovwMxiITRnL2/SlDpdrOnor2GZ1XagIv2YqdE
L48SkBcbj7/UhwFLXzO/usa7uYsQHcC9gqJiFu88S6YunwxVqpJcASBzrhFUYS0OoR+D/ZjyOLCU
6+InSg9WDNScBoR6/+zLWyIm8kC+6GOfg7XOz/m3aqFNGaMdL+YBwChFzULFdZwafGe/gndnOKGH
F4MJHT7WnSqEZy23179SoQ1d0z+oVVTKTGPIIimqVEfTk67gOSOyLfc2vWae1cGXgwy+ie4nLare
T8SNGeh0e0WvC7eGA9ZVMsMSTjWA0cF6cvK9zLxOH4giiv5rnCJ+oZfqOwd0AYj7thA2gVe5Zlf9
+Iaca0YFNj364VT/vJieFonB0vZP/fw+Uut3qZM+fv1WR1z7nfqVx9gs2QYaO9e6f+BhUGlcQ0c9
sYnlLDqC5z4PG+xtRwl9voSeZI23TebQls92FaBto8A8g3oXrjzuf6KSagLchlJcI/jWZb7YNi48
OhSKdkVyckQZVWhVFPdugoRDuS0TjuN6Tgy7yEbM1FjhsNz8FtnissqHwmljO3ffIxYwpHnQHgFN
8OsTngoJ7XN4EDWWZON7Gxo/iRefP+7Cqw6d+7vQYSMprDUntm7jYnHq2rbHd6xNyMeWmepZc3qo
qzsKErxw+G2Yd1YvL8K/SgW0b9Nw66paW8c58UcV4avhIUG8Mn1JhagpTLSGUgWfkEpcK72CCriy
nlKZER3DjL/OvEvNxOjeZR5sP5lCa/UipesnU1q13sKe/GLDvZOBSYPJqKXnBUTTEcZmyL+aXYji
PBulL2ueBV1+OmRwB/z5JfxDtVNPAvIVnmt/Qg9y6Cbnvnd5tX/1x599ZILK7FGoaF9hwQOozxnI
fTJeh6Uwl+bVX7Oxh5wTaOk29fibsaCAIOgefZfkaGuBpapGmZMdJMj30xhvEzSUjFH8eVUmEQ9A
QOhd6hOEU2A4HsFSSJqdGh/GFAo3zfjnuUxYh0lC5d8Ug16U0UgpICOHXHGHIg1wLS6MjW1PoXWf
e4GNmkOqDMCeH1xx1E8QPYXzXcz0R1RPTujEJ8b/s1N90tQHCvJrx0Iyis8l4wsyX5qetZC75uSr
N+32bo3oDLuQY2DlnHSvcq57OqGOHwAm7JkJVJIP/HPYyFIa7DKfwrWU5bTmhIO2XVXOlRQTGcRy
jVZiJRq0LgcIfae0tJA3eJARZnShncpqZU4FRnWWfhWrnBppNJn/6AZfh56lXoEfnRHkXbDA8DL3
9InIqQDCm5iKg4EYUeYrz+hqjb9Vph61SHgertjqsFP7llOooZC5nQYpTfajHc3WAC0Lc/CeOlWC
8CRtMJ2uWTW9il8JbC6kB54QEK7R95fYPFME3JbPGIo3dsP22fuElgd+f3hvCcBzzuXvbVWuaWUx
PUaLIG0zBPLRJ2kksX7aGt2Cp18tLFjUd/0rzwH01aEQiUQO9yfw7WUrs6tXWps5q0O3lxAw9Zjw
qFos3AAZCIxja0X3dSUWZtvrPESnw2fyzqCgBx1wTVGPh/Qz76Q+3l8JiPuvKXjG8odhNTjLsU9m
Ju13Oj+Dq1w6W9PoaJzym6WKIgbAPeXi1cxhvBy3LIiuq2muZTrBEq8xOaTOAk/syYY+RwxNi91C
dON0KWirHfM90SxgRDBMpqJFJ/yV3I3MP72xId6aafuBOOEflzZMijZGO+MRzvOQYX7eT7VjTMV5
yhqeq35aENxMq92IcCg01xybjYtjQ7JKmmBvEI1yhCkIbpLd3xvDWydYwD3Xg8kc82HysRcygOnu
bS74lULcyKbka3LCawyDFEzoLudlCr8N3oJkIg0H0W5Ydl/2vT1c1HKCBfz122sYdIsA8DoA1UKB
+C3RhH15qufIqG5mYb1xLB2ikZKtL0vBTrZ4tMlM1bvl4PO7tK9j0hVbG1eSmamDo4jskuz1UB/6
56OcV/2vlztWkQWIzUF1GxfSNqiEWtrW1Xqe+o4R/zOuG1m479+TrDozBh+P87VoHod6uELct0dE
LhlFiSnpK6VgFaLqKWLx6S/OcP8bVKrhDfTQpgdx2HPs+/av8BktDHRl2eo7WpIvpubJrpo5PuhC
/m8AmkkAk+N9PM86GV70umQP0NN6AXA983RxGB6qzr1MwVD8FGzFU2+b6xkhDeF4azB0IHbkeci6
RqgzUXtZz4XSx4JvmV6NTAzXey6nmr/u9oOYHBOoDmNDWHKd5xk/twGn/P4fznPIhE4y0fpjBIX2
XefrfcY5W+6VZRkHMkPFHtDqsK9JQqBPGPYpMvxGm+BIqsr0xc2lhjYv0mln08V1+dBLMwGiirS+
U1pSQWcXciBQuaOjCBBPvr/mJxT3EOjWIBDWx3fWjfxEqYGE8GINZaGZexIt1kpt+sCMVO5XiJ8n
kozXvH7jLHmYh8/aTpSXynP/RBva4ggLh9difQQncYPE9pHbSlNOVzi+zKFbE1NPCfZB2vdhM3NQ
2tV/hfaf5wj86T75tqXTRG2QJeyN4ef71hBGBPqtp5bp7nW7vvQxPzipVLfdifgaBwHBgMk0nox0
7h1LlzMkdHfyuJa4R9R+WVHG39q9RFr5hybfPfXBk8ghMx4MdJkAQaFuWLPxwNqmIrAaCDJBB4/J
c+lKWcIDEG0Xg0V3z+Q5y7sfDeI0Sm2LOOe0sZ8FAihTXEi3mWiOidoUsoJGA7OFHBIwIvGkUysI
OIEtmi24k6ubH5iEZzpXQ6UIPoXWQNvpyR+j+rAe9uy1r9calapS4N9cE2oUnrCLE6rS+SztffcR
n7J92ndhBluevACOVXvD83vcDXzseTZfvwxay/7gyQM/qVv/rjz7Z9fRJrQuPwZuovsIoZv+bNb1
7dNs/e0wsIgAXIssS2+xcXuLozHoA7JqC4SE+wOtnVhFOQqvyUhNKaTHueOX0XNTYM8v8XNIFktE
3cYS3/G/AUTICx2KhvQWrK/W5otYzfFASrjMn8z550W9w2P4czI0t/Qubo+I30NkYjIc2t9yVkaZ
ehq/nTIxsESf/1CV9mjNqizEUuyL1CBqDQ6gUnWi7zn/bzubH80qPQKNcWrH/ygp6jZ7ZJb5whGh
C65BymIYnix0OwbQXJin4o/vh0ii4BFAHRKHz/R3FteIOOZ8L/Sp0bmuOa4xJe1aZoOZcKjUeatI
pzptlywmf1RkJQnKunjTZf6MgR6cEPzi9yBX9nKqAoLlEo3tSo9FHFZTPUVgD1FvdAb+eGmPxSKf
p870f44OTqwjb1c0XeLbwKqFqXa7WjtPexfm6P2g17jhbhgggo2jDJA4Ztz5ZCwOaeFtuPWeb7Fe
A5AHA7fKJv81HEGXstf8dVXqt46J4snAZ0vUL69+/jj14uHijTt5jASQWHjLRaceTzkJ86lNIEPg
tXo3x0htpRUM1JxwiRwxt/rOzICbwNuQJPC58HN1mOEmzQLmmQ1Y2f0q6LmU41dOUCNo239Ferth
lsXh54vwhGHlhLS13bCVxR3N0Eq87zWW8Rl9CBLuws4vT9ONT2oJH4UmZTixg9ndOh8rdAQZQ419
1snNi6GMwL0x3xsP6MBMdQwFzD6EDP5z6McoPY3it6UVhRuPA1Vt0uXoTfX6fp/n/2HpeyI+sHU4
Zan8pXcspbNI5vI/BKa3ccbu3Xv5UO/EVbjqIXQXJoykRz2E5agXUksGlFcLonQ6HCC2i7+pYHOq
xVEtiJaRnNisIZdnFA1Vg0L1ccWL7wmRMeiHtK09ivcgonTxl7xt7l2Habn66QCbD/YwpNHNyArS
2Z433enSiakLTeEJTUMIfQb94t2YVAtwXi0bliTvfRKlgxv1L9C6bkxdbQggjwnSOh9ycRK1PHsI
htN+JOdnxkZabrOUTiecgE/yL6heOZuMlw6E0c5cKhWPL9XlPzC2O1sgAwq+nxXmqAbySSH7pD3+
SB1uAsGnsFeRG9u5grbCymbZ0gOt7xqf/3bXVXPAv52k3PN5tDuhWn3d1DCqQ53cer1Zw2Pic5GV
flNAgA5Z0jrIgn4DWITZYisql/LcYI4dapGqSYRzB2tVq7inQYjR10FQkybQjHCbvbRwpMemyMM/
KzqdCjO6Y6bYlyYwixI2kcq6e60Lt2jMDJidWqPiTbxjmb/fU8xXKblosb21FsDf23XGSfLZoUup
tm1SXcF1u33bN45vsA1Mg06K3Xk/W2XxiUk5D9Xt1qZEftJa65NslU696LoeWubn+hkrYSYoXj8y
fJITMUBstGMVIlxClQfKw6B6xfhwrcBvmXYAkHJ5Z7b6OB9UpHISOyl5EPTwB6u5gjUiQQPVAPQz
W4JA96LXmysKJsnTn+c03Yes7OJplBil/6iHsY5vZggmfONkXkhsTc7vZdgGHecIBhAyZMZtVIoK
YHGcuc2tgn182cfxX11m6f7MLw8TGBF5etU56+ZTnLfXREoZeEdNAu57Y+nnCTdTX9JaDHKJZNQj
PTeV74C41m6Tyn/LkPelKNszoGr/Iyeinp79UTQzDmC9jD52xEUolhM9NGeh0TRXelQ/5yahOCmj
RtUSzTRjXEGC9WuchLghAnqN+yAyCPTKQYX9xhCLEjgQOZAojsWr8c1VGWWGFZ7SQoU/B96LYYRD
npPMQ2vbc5ef+HO7UBEqbBGNMtFKZEu4SQ4y2WBy34AGPRgLqEHNut0wYaOgnySTvRRuUa0+Vwvr
/gqmeI4cRsHDjGWqzFJwJrPCuGxQKlDcHCtcirrK0NFb53fqghsdr19+zMYRl6dai4lHtly1S4yP
Oaw8aiW0hwRa/HKH2JJtzbMUKoZ9FCF2xIbd/Hc43bnwTowonLXAg4IHb9bhmh6be0umpsl7Hzol
sbS8vU3sC2usG7wr3iIZuvmRUMP9Ip44GOYRIxs8okQZVldwUhwQVBQqLao2ZLNzKceGWdZk5VxK
YxxVrapafBBDpRS/Sv9Xdk3+epH3omhk0MWiiiV5lr3T9+Csd9iIKvwMCHLYLwu56Rf+oeajyzf/
Nm2oZ8qQQ8TP8bRd8w+BYp2FYoIiN3zBIdqV/EvxQo1EQqsMdyJXVwjufYzknyn5a+ZlFsK/uxOq
AB3ro45PtDV/Wf2NuhsLp4RmAtoxeMqt0zF/ohFyYSAv5ToA51UZy1SGQCu8iT2ieHMVV6C01+Tj
a5Be5VkvYUwkvkkNVxCTY+cLQ4X4oEGn9bMrc1ryDKaG2tm8v40Q1beAWFRsa3ZuU71xipXbnGVh
oZlnXQfCHa+Dw8giSVswpj/01FenOqyY8AGhwsBDO1r//pFB0VEBuXSh+JPaStruYxkvrFM9J35j
2yF21CZJJpqnfMaf3IQZNFPLzO2iYDHsBAEGDnNJ3By5vvw0eNHqRrPoWvZUIdJV0c73YK0a307H
jq7Jbkr10yhoJPgHMPrsiPdleOSwGPnHnoB0ag6OFOowYOEqBBm/YiFnxaFx5fd+VdEkrsDebh/j
XHrIdw8yepRhREn1BwEXKad1hZzq+YxsmoN6o5N7+YafW3KcMOz9jk2igmPbeB3UlzAghYwcQIWK
Ivo9lDXRCQzJVkmFWSMz8GHLRuhexlZG0WMPwN7m6K6agKNmxCXbvBuKPjyOcKpIW+Z4JKBzVTzH
H3BwX+vzZB8sJQ+psNDbEHG5XOpBc2TgxmJSUQGYRfkBYoBZKYF2oLdPaBGQ69NMVMmNi1gO0ChR
ZVM0OxlTPo9Ts0oG1BGl+hni+AfmRaq1M4qhVluNdFQzBJ4FNjP1HKL6gBntmRwFd1amvOKJ+G0v
H8Q6jY8dyT10wTChhU5EKV8LPZ4wVBqPGWaxkM/99BfTBK6vQ3pMq76XXeKMYgtPaBYzcOp9N5+X
WPAo4wvOibayAkRqV9mFvERne5Vc0+3di2SiwI3JeazjdWNAwaDG64YSb7gXN3TdLPH6K5q7bUsz
aDeeIEm9djPkb5FqS8I8el0zBarXwEo9ya0+vq1G5AGGLufHFvpi4ejMlCQ5YiahurRqfXvR1wGh
sr5r8FU1C5myKf/hFjzaHftz8lez9txqwd6PoFgG23LFy51138NKnPBHdolwJ4lfv1DHVafnn0MH
QzV3oAkXcI4V8C1dmsv6pNoLfW4bYa/gtmFkbL937bpAGzX8BE6VURV8LTCPXW1CzTKtvaLS4MFl
FaJaVO9fPvFnZ9nVW7Uk30dYt/MRmtfj2bj9w973+GmFnBmbPbD52nPVQeH729cDssV4+ZcJSxP1
z99xwX3LuLiLGfT+onxs3FlPPcKXRDdBWbOqTIEeWvpTt8WWC4Rj0LIfsgon+lYrLg+KNhO5I7mP
3DqC74SKGFVfczuwGp+gaNHKIGwIxj4Lnm6731V/LIySAdU5C+SOIP2EUQIeOyUTNJuS3GcCUpIm
a5udaZVYCuCIJ48t0YXCLaqeCC4SjjzEGfDrpVnftlWQiHxscBWM7PdkLoN8LH+Zdzhgvc0TVFaS
q1LLND+d2RNNMvAAAhAoeanN4uPiP/DFRcDXv+YIW4c7tPPP3/vY+R+G0kuSKo3SIdIXQUy0y5Pp
AMGsL5b1Hmn/IPPITpz/nPcR+Y58UeLLaBYeUmvrv5ktgd/f5Wce9pNSIZgT/rLPzZVrwQ2m4HDW
6S0yfoNKmpXhZttjyBCWYOl/kLXkXAkTumbeNN/IKAoHsTe5NFv7dFRZVyoQn129NaXj87roa/6S
6QWeg37kjPsvg/SIXULzJLNtfROWp/IXkgwIdKRZmYYNwZA2TQWI6GJ5aLaDW2eC+eokdXhUaaW6
akeFn6OUJfqU7RBtvGGy+ari/8uX3Mq2j+WEOi1iCyb6oxzGq143SO+00Sff9nKtAcqqTAPoDQzG
1ZYofpPSYqKGUiOuOSZFZgZX0ZWtWFp4D548Orh6EmZV63NEjES3xrYC4mlySGFrX+XuSIxEhWiT
smRDlRPYoAZ/8uGmmKWLRxW2j3xnB8jXOgPmO2PT291MfcCRLwp7zPlbky585eHXpP1n0ULyim/6
OinymqVRkDcvqogHxtAZcHLNVyu5CY9843usF7S9uPyzFvFLkC1GswB3Sjld61rh7wi++5isxP0B
uRF47IJJ5yDncIR1WoxJYQpMwyI/xurORKYRju1PazGO5sg/BnjvHbFK8HTbFaZD2LzVbatvQsw6
wOSaWKT6xlJxZsCkrtbkDdRlblAjG0lEEMHyxLotDDw4EbVu9Ow3FUIRGF9Bs9c5fvcu/ZVO6gDa
9Pq8xYIV1rOD8lN9nBj4JCBOSdeUWoeoL8nBy/shnaWAZJo5FXTewG0ERs85SCPXhiF+49Oz7KNO
0MaprkVLtdgZlG1WTGiRvB6YnPtz+bPY9teOMl9EmHeufdGioijkEhIPTbecPIhEZDy8DPnoWtId
vY9jC0x/aizTOvXVL2zL01C64VpbqV5VPR3iVKnZpVU8jMVoZa0JKnpwuV+0B5ELFQdvHhPgf6P9
Qi0XaGvx8deALGzL1B14lvoi0nRRzb4yMWEfk1wBLhOvMvqY5jtrpU6LOvNPHfz8Qzj2O5CtpMT0
AbMTDG2YgTEbRLLiIw3JQQotJFWKgsiRQiodsw7fUe+rbTjOD62WZVLPZkoj2e9RMdZ0Kbbt7Y/x
9RyJ8ozguZ1rgmygOWCbbP7LtuA6JrbyfHscMGPw8Lwj+g+n3XGVg+EoBsf+kvLEbQIswLqSB8KQ
morO7g0AqQnMecqIlzu92/T9YkXfJPS3N6w7HBSGSuTBSyCBjjx8wjR2Mrvcme8ttrFWFS57XR3y
TJ3SZpgWpEtVeJTIAXKwesPQX1qjyAAhLFqllmQ1jlVsA2swcleta6Lh/GdcoAhNDF2SfvN6kVcy
tb3ATnI7wx1AxQgIlttJRVilT1sYNgrR8wLDFySLkiEbLbUQbuvbYksdkCqclIxqRtHhfNTyS2vQ
OdsP+CWrWrgWH3xl0Jaz//FbckWyXFWQ5T8zCVP59vRgaCv6v1WP9c+00GlsrSbFdGdIOW1Ewic0
5TYdfKPJYW3d7ODMKp1SUSnDIK3Qy/v1c2sLYSGyPULQblxJN2DtarWWLyx/DbAhpOIKByo3Plni
fB1+tsV8hz13LZzYnZEpX1jLbr5093lGkjlDE9GOadomi0iQXJfHa0H+smI2a+uJUh28lF8XSRsO
LkX2rFyFozomor9bStwdYB4cATUB9Zik4dkrYfEEPFDn9KGVGq1yD9uTDO4TYLqQJUtF1lkwrR7I
ArHP8Dm2DsgwyYptBYGBR5V2Y3df53euC1bd4sdc5rZ22dYVdQFo4LKsF7/hAQjYeEBIuX2ua1jl
D2LVuDcVUbsOKVZ7rkU9JNEgxPRUYiyAI1vI91Zm6I2abbC5lkXtgkPgoaAGs7X/LgD2tAScOQTE
Djj4gCY88ta4DTqG+sxoSqTW/wdBxicr9hzcNIV0eOhmh9nRrTmci7haX8LMkF3edDxPLZtGBaeL
KuP0GFoCXsyvVxOSWQXiMmKibdM5qZXNroZfMXr9LsUb/k5HL/ctld1BT1zPys6RYwwXdccHOgCg
tnpBWcqmIOZDVMEEazwvu214qmWFHZlM6oK8QRS+qs3V5HMeKLP/LB7JNFvpSUe5QKA6em6/0NZi
nrL1Djwik/XzYhNrIDQ1GVQ1G7sZ4mY4NXshoAjMQNN2eZfB7Zxa/vqos9K6Qc7lkUViBzGLx/u+
JUVhfnz0wc34cflavgxoAvsZYUKooNyGuqwHA9tqs1YbvCZTaiXoefY0vIFqu7zL4oEthYxMp/JK
1mcs+ojdOI55eaWyqe1+Ya//HI412opH3RtkcCzQ+De39H1Zoq7jtFANw7DZXDcMG9Kgd+mm1wtX
/8fikq0/4o1u2FtzOIjrKPcV+PqAoRVNCfimSw3ZRMngLFLDRVuXtmN4TKeHabpD0UDdiKKIK9wv
sCR9GK6TM6UTIM7DAv3LHZn3ItBN62v+k5UBHF8tvkF1065az1K228BxGEmlm/miZLSw4rVP8ZJ+
9ZLRzIY1ksgmAVx/Xo8L/LChGlnTaelleKbUJE0l14VK3Bv8Lm22/J2fvOaD6STX7q59xqQAFemt
18Ttv+yB/oZYLqPVRa0nQUPHpEknlbX9swkGaFcJJ33u4MWOWyQ12V5wyH3/2J7Yce2xYTSf7s8Z
pCSNXz0yTnN4TeGiqHTPxJ3fcFpGVDavVYYJDnvILqrwh5djQZRxty+6q2xq27eUePg0ZlqzTiuM
jzyRtylne9fbYpUEgv1FiEugSodLnXtN8p7WmP/ykAs9XXH1vXKUW5IwspXCUettUK72fEAfZ7d9
gEKre7A0XK20kW53Js0XoYHRZaZ4S0G5/+kU6dufifaqXhKpB0KlEKd+f57s+VW09AM6gIIuB/p/
/P3Hdl5S6M0sdxkJbT4kw5RdzrQjxZmpcE/SzSPiMzu8KYP3Bt9Q05hUqDEj+KstS1jJS6w4zrlC
lRONtKJqdUHf9j/BoRaJ9KU1S41RYuQNX8cBdfT5O7633QiNgkl9bLUOfIvcZQ6x3SB6ER+8/TbM
hMJjOY8BBTDWA3xtkXL5R3gGTaHmpRSm6dQ6R6Q/QQZcOdO43wnjyBNLRDBmIoTwDi7UpwbncYHk
kRA5s4zTI6xYQdm4s8sNpDJQEElgstIki98c9r37yYsG/gcEuT2XlGAA57gjc2ayjFJWBDV52ZBr
jv8CB/5UvNnJ09n/uXKFuEppxZVKE+MdGNUR4lpgnPFF7dAn+Wu4DV0jS0Cmkqf9wfvJgj06SaW2
cfxh1CN00XAMnKyQ+NqetWZrnTy7zASMRVvgICo0ltVP61F83VZ23bY9D6PmtDR/TE8i0NEf+4JR
tjliPEwYkFid9iK8OrWDlgb4JxDddPxT7u6lOq6nNJydesSlFL2zECgNUqkqFkA92GEjZgSNdg3X
HpCWks7CGQR0lkmxWITNhCmcEWJlxhgN3XzoUHjpJP35anO/GOmEaeDW5l0rfAT4TqBCw+uhrm/A
15f4QUB3UcsR3zdSxNvB9ZQBBaOvzRk6/YgSsTkzG2b4Ptl2bBp7HtgIjghCK0CMuil7aFHdbhm/
GqeLX2u7GjjiXz5scm+lDUoRrDTSfoHhTVPkJgLSjXVIYo961vQXU4gwMG6qpEWyw+IQaPAbfxGV
qVxJPrBYvv2Yfa7CtUCuL0dO4sd6Mxyjxvs5vlPP5hgeRUVgTMZ6Ebfw/mSgv4DmdEkQ4xyttiHf
NdJKUFtl29XKygbepz5C1xtzV2bffeFHxpV1DP0cNmwF2u2biFWF5C3tQjqlcv/9aVA4GreaLkgM
06uNsHE+7QTiqjMMjp1c9LT3885VNok62/+vDtp6vIyqGk8/qlFkVki4OUdS4PU3BKRRk0nCCMSs
M75JyI6g+5kvrWeny/4DUTPjJEnBP2/dyY+HzAvcd+k2rIMz1d6qEHfOUkgI01DMP7Ne0s0sxM7b
EmtaCrq8PjKTSNcY1DL0aLdew2r+SorQgEcsJw1kCizvBIWeO25trhJW4l8rU25Bm8hJ7JjJWP/O
B5uT18BA3hhsNpFGGM0MjZMlRJHI4yaUjEf6c6lCWUcm4k9ga1tGltoeq3V1r+0ZVXcOmaLCFPJO
hbcsSOtHt46rsaaLUnGkWfOMdgdtpJjwAgezSRCe4AAw51bWQKfNgQlD1JZ6lz9AT4lJrJBotWHW
/gfuyQ/V9J+EsIQUr+iGYTn2GyxuX2FAOINlt+TJFWHdHSklSOPIkMPNEBfUw5fD56x0//i8zSIM
PQ6eF6ld99OTLBHCtzt/U8WdZEixa2JBgRmJF0ZCXLbNEVMoJvSaeq4T3QaN8CE/fza79KkPhrZr
j6RlYdi2XxH9Lxf2fVdUZjjalgt87G9cKViGwk6ZDbV1YfPeBX907+TFtks7C5KLyXs3YIjVgbMj
CoX2578KZsP4sAwv8DFB/3cW773v9/ANCt/2YnIVUq7YbH5KUvmZslqxCDrg2SCQId47AkU2vNhD
iS9Qdm1SnX8sknPcEd41rtcNE8yQl0gOtMCxjLIlVbJlALyKB2PKXJZpXyLDSTqhHv8J1rNvnNPG
AHjolWtazRfWknxfBKB7l0JbGVI3KsAtnHc33WQUOnt9q35QgXk4nqH0HVj4o+WexqoLFGsyHPnE
CoC1gyyPdqaPV+p/zK33ps7wnyPW6JfLx0DH8gWRG/Jxmj0OK3D1zM+FKTf0zM10xegdQEc2Rw6x
4vAaTOcAIASp2qCtKEWjqDcL7RJE6dumpYggwRLyG95JogWadF71Uwzzke3FMUS/I3vUk2KHzSvd
5b1UUHx39ZAusI2QCglNJWqOx54iEPaRwS+GmTwCLuJ4KFE9sTgcyIPDauxBz5/XAvWT1FbfvJz3
+ABHnso1BKVrWFdXr40JZ770Z9qhiCF10CWjiYfXJf6kOkAJzIjoP+Pv9qja5f1RYgdsPLoim3OA
jMSx0NNQCb1YONQaUZEQLa/tHhlYEkhexoCVvRvl/AdWk7cOS1NYAq17PA2fqu55fD4DEmxkkFup
Z0Kz+T3tm6kJgbfkiDBx3M76nDYhfhzOlGHF6PCUrUPb4aTeYTt4WVzwMGOlv/PfueL/5NZVZdm/
6ZjOhhukM3wNmzWpmiGe/cDxh9V3py7dtED8DpvGXMWuAi08/741JT+nBAVYzExNvdJPTVVODkKC
Glr7piX8NpA6wuURLEhggTfBZlwQ0qlkM9j6+GuXbEEeaivCjBe4slqjf45t7H5cGo9wbGEBDk9+
AHbrZ0PU19bPpg9+XAoekF632KezFcLQldl/MCcCwizL5MAe2Ko5uTvyvsnynNKuZRVPrgJ57QHL
oLjtOoob7sb8Wc1I9NRhloZpfd9K85Ni94cB//a0tK6KoqhgIl7Bd+t9gi8GNip1FfBzlGf3F9sr
2quZu0+NXOJFXcJEjFhoH7nIUFH5RxL6UgCetr6fGBqDQCvcW+BEiyVXrfbZrvDfBk1CkXthqp0a
X/jej7/RMjrIdb+yAYbu1BWb882hzvumOFqv0y33AXX2c42WorqKXR1zxnV2TNwab/c268uoBN+g
hv9gUxYRWmrM5WwQ4Gt8B87DBnPHa9moVYO1ektflF3ZOV4LUSIo7dWfZDYQOarTIaSLsQqDAfmN
QwaEVAFOO54dSjlmKi83hKNgRDt6ydsrCeh+YCosV/4UjAFu8Brr8HJlG6jwl4ifDL/Cu7p3Tx/Q
RnWBuqyjPswcD6GKBdrKEnMRJ2soH0t60Ev+xRjkP1NHr8vXoG9u6zYcdFN8AdhNpV4oNZxFF1in
PN26bm3ZMmTAxtCbXtLff0n0evdRNk/H6vABHvhx8d3pnhJNMX+S2XoqeamqXkxB5mhhDLHvT27R
h6NEjie/Ekm2ijSQkh2HRuHln2xkztTTiuTzFjtl4zY3FpKIDiuT8ARjjlQDjWyoEdTJW3nd/Sk6
zgL5SPMz+clVURw/YGZL8ZY3bwp3EaWrBqd00PSxm1qftcSjjyzFwsixlvcsCdUwIhr06S6d8vxC
5YLFuyeSpJHqelyfQj+N7c36mvMtU74Y3oZNT0HHdovuXJIOhXaX9HvV9lSnpoL86jhM/OmlDQZ3
GhXhIe9/JWVOI8jmA0c0a3BLuPutRNLMJ7vvdihYyJWfhJ5iVUX8dcno1eH0YetrcNI4Yw0JwBoi
Xlj92CDoCD1GXT+1sEKihEJlp6Lr59p1HrguqgDH+JuIVTynFDl+vRcDd+s/OSXDYcUvlupqwKoR
PNT1qE2a9Yh/nu4P5FJyfG9+X6fKMqKzWPoEYPN8lHOICT3lgah0Krw6y/Ymc+lUxqBCibL26QY2
95K2dwUw39+HKK5X8kiOLECFSeWVqNGB1JZuBP44fZ9wHn4CPvWOkQcaO1X2uet1jF4UbtIr0h9o
W0YydS9w+xuqnm3zsDcjlKQE2j/MrUo5HEhXAJk2vg1yMXvR7BsbKzSKE+92Kgnx+u94CeVl/U5C
bU3dLUWO1tLUyIAWgTxGsj8kPNdeqI3hOh+hnWluPUeFbz89Kqub1nHElNy18zYTM9sQTzUjLKd9
c1xagT1Y7O2DpTDX6tN9Z3K5gMB9yJoVgZ1WyKaFzhnt5cvinBuqyKBHRAeCLkkV/BQBkzr3eFno
VXwVl1Tbmn5Kzq/v5orcne+/0Y81GagLK21APuLHAb5YwYpRxCo1H/2Fy+RgdQkoZbHff2oTKXbz
LSb7BYxJv2wgpsyVciZRGIY/HDFgsxT5UC+gG3isrJmXJHiNGBOJC6hU6+iRr0LMbNmhGn1D2o+I
0tuRUFcpwlkCFRIkI7MRIH6aw80te1dVOiXImZ8mFPFvS+CxiQhSfmAGgV+GkO+75dxPQeM6JToo
Kv8QGw41ve3/niQ7Wj/U0ev94SBrC+oN8DA4f1PASrxOcfRGnsQ7Txoaz/vs8raEKdZm1Yp2/k4N
zf0zhNExBADp77RH/gymPgvOdT+ZiDpXNVwgvf0lmqgDiO/Q6bxqaeGwwU5qxtr19VuJEinwO0ne
Z51tPwAuJZE2uFfnKA3KeNad65LBnS4KUuZBiKzi2PijPha014HTtAw99HU+04F9zRKfiHLkOtpJ
rcJ0zBTZRh/UzV2U5Hx2ZhMPt5w7/UNpib/O5SZxi1OaZMGICw/GWpvKBsxwgFd809KA00VBv8US
4ZfjqS3Fa+675fLp0O6yczDK9APEg+5G+lsKandJLP/gDPi9BIT4ZQYqQcyjF/+VwWExs8L1QZpi
wHCf7KNE3jPGU7ldzj3CiRuqb5jQciIb77AHcg8v8+4kLSZGN0KbuMW1I+qW1Wf1exIdVTWJZg28
Y9eHdHJArLikP0WJ3/s8m+LcxwD+Nrc4uYL7GfKhRPVZOGitRegcmw/D+mbpcm86gYv4q9P9F40q
diumZ2djVkqTI2XiVsblwgXbcxhpwab0UeuATmmXSm4f7PGoYyKlgAE7CmmBA4Sz5rdJCQoNKjC4
yuUGSajFwrIB3EJIReGkvXAuRYFfpglBbzvWgIbbzpgBjAA52YvVU6pThsVJ9ULAfGSWANj61CHd
Tz5Vu3lAyfM4bIJal57sC6++dX75oQU3D+jz902RdDj7wLu5u3izZ/mHVgrvkuVyPZFfg/bOAKjy
BeIHd3rNpO3ZG44AEV86QlOy2b/bOSZmiNz1CfEr8yt6GjHVw8h/IoGqFPwwWBqX0q5eMEa13ZHY
mvRxXHmn702HpnBqj/IiV28Esmmy+MaQPSVwDdVYQZHqg7nW6IDvQhIqNuZu85ah0XKMn0mufBmm
NEvCNxr6liZag1zXs4bO0D4y3IQoLOlF8cus/Fc7uGMyLCxUvYbIGtTltsCVstjd62v6HklYGTgY
Ybth9VnaUevY1rPAZnZkiCR6iMkS4g84z1TM6fhPTEhM7NWAkp5NCWuvHCl4ioKiPVtnF5NokwLI
T3LcxxjsPY3blK7dK4k6fsz49wN0wkYTyGeeb7yB86EYH9m38RgUcPeeUghRq1fdbe/E+MrC0y/X
DATyXFkErk/iew1urXMqJBTrlA/jizC/GsdugqZkByMzzTP7MwNwU8VsglrFWIDm14jDq72HD+gI
QFLt2tfva3NWzlj+UfLxuqmxctrbHxxuv72zjKQ0cXnIpkbYNg1a7vceF3JG1P5uasHS4rpyqNHa
CU2+YYywxsL2Z7tpTZ2KmgPPh0OmNV7AzGRSebVZc3m/GLkJ3excKpY8L2MfqFqkGxNlhGnRbml0
ZSacgzn9wk2BIXz1U3nZx9TftLbN9fkw2f3b5FwjceM2H3DY01Bu+s/0ZtyYH9HjMkq2igCBjjqh
BMBz5Kg25ZDnjXjNL9wMTK/YrJvwdQzYWvpV2T+W9FtAi1agx1eUcwbwhp9x2/2RfZDRlZffXrrs
zctHvkg2q5Zat/siUJ2UyLnDii3xPKgwNRKV0RlHnXMjR8W2TCHNS6gut4vrx76bOzpZDfZTy4iw
UXB2nlI/yEHcs2sWvjcgWvf+qylpcPX7QmYpSXfd+Nao9Ji7Eiz5jiHNZMkhRcAxhlN5Jft/Nh22
iTezdJT9g5TRbQSI+glv+QELYKZIel0vBZCFWTIPnZCRolEE18BbCNzM4WkzLc51ESl07LuF5PrU
iyYmxW5GoLnVuqh/KtNML3fWoLkRXLsq1PYI7yOirJqfVEqkvIM/zHtQpouZx7WAdWhIaC4/1jzi
8YtYDK2qy4jiM19ADi9CV3+eukLkMRPzjV/JIIY6rx2wzZ2NgLmvYT1Uk9GVZ+MQoTVfIQtJ5i/S
dbTP1Z+j/eT6M7tonLgDfqtCiiNo9yHDySLinh5rHosOPnvVpBmvKKijtor+YffHunF5Rpc3tQGi
HjEBlU4ZwPmIquuBujt5xL5fhyzDjHN/nmKXDZ/s5+ZM6RnBHuMyGQPfvc4YC19TgtYklv/5/GHC
d+WA4RRIeNDXhbP1qpUfsT+UM724ABaOAfRV0WLRzEpsOGVFHfpibslXkk8dFJurxVnlYx3te9c3
zijdPmHclfjKWrTncHCC19i7RSFdSufaww1gizRDdAsnsy5juS2N1Bu/4C1RSi9ZL2u6F20mLD5j
4YMluc6sC8DhPnNZhYkzBdU6PwFTbot+GMRYc2GmNrTGkFNFuGpUkZR5/8yJHVOtXFhNWWOZvibt
WHgSMRVJ/hJLD263C0xPccS5q6yL4bBjxJ367O8exME1Ix2fqOGvzy9YHOPgqf5Gkkb6UBx8tGUj
SrtmT2hlcTYuUPdNb8vqjqa0FL9q9Ax+7/IJXbsDIUv/+AbNEUSb35QbaUNLg3q6XJFt0rav5j43
1I3QpGTMtEKWl86P4I5urQp5FGKvYHanuxXVr3OVE8bn6YM9UH/VW6whInmzQMvQvKOVA4Z56UU5
EU1p3qwtQVZ79QN8DAgK4ge3mjP3JAEbnzFuNPGgaYaHQlJeTO2CXFfNYrDt7A5iqHRIEPWcR3lP
w1ZdaCfWkGoFNPH90SU6HtjZNAbxlOVrfY6P03DwLdMSxa1nofrU6Xi9CGAz6mf7TSYhic1Z1Te5
hfMLIWJH8S2pGT0TTynkVxBUiw3mUBDUgsIgthRSuxhBufZngZtaNt8nxKp/MSMipWj1QTs1QDaO
4PwwhKc54bVRq47yzNuX1x2AxdRyjlZwj3nVmZ0UWyu4E8vwlyB8ZTOlD149KI+iYreFZF0OEZTZ
s2z8Q1sQAna0cNpB1Le7BXWfgf9dSFgyryQ4uUOTRnYikyxfdaZ4cI7bIJ1Dh22Lmspp2j7N1jKn
mBk3tGHEpY2Ef40w4Uvg/OD7+Izn1EKQ70Cmrdn5u4pIVdKpuDY/AR+2EV3i9Z07i39lMu05XB5/
FmAUP+Ar58yZOIgMU0XPctzt4Nc+sIcfr5tI12EnCveqQ7DA0Pcs1AIYMvYVVg4imdMSAxhjE8ev
6+I5FOjvMkWIITE+qnan9Gg3+JJpw4+y+4ZzQTs/qd+Iqu8JGBqYxY/3uOLtYkJKJWwLcPdKCUl7
aIvz0R1bb6Ioaw2hYLm1WHxLQRMQ7pkLJeBJf4IA5HnFbnEjlxw+IlCMt8GALChEbuIIwF30OJZL
gurQO8PqcpJjQ3tDQi66E5fLmI+lMpP8mrNzc6noU86rxcmDdAf9qLhIPpaHXRIkoeNllTgqmJsy
cBgvBk4bWW5AAmYu1NoeaiOzC1J+gybZbT/BIOOAw5zzobjhro83yR3iytnxOj/tvbQDOpwzjrdQ
VcgEl1lN9kfr+hyF27X/4x+dqhDd+bx0oJ5z8lpgaXwEJu3MOXL2epvRdmN3cnkhgZQVQ3WzYx20
Ms6hpEnMON4UfRX0eG1LYnsdiaveL6AgBaFfmjiRrJkEHG8qy/5u6KkarLgGkNf8RhXwRU3QSJ8C
KoZ5/n3ZfuYk/5ZIgYn2O5Qpigs4focGOULKUjW3wFo+aI1xQPl+KNaiYG/1qslVGEg2wx5D9DNf
KQHn8wnNxkqtgIwtAOuNtYp3/La8l4vhz5wVnbnuLTWrjklYckNhCXylwEb4jtXvr5LAIlEmBKSS
fdQDudcE8OXRXkl5Hk4zyIK0e/3L1zqhqYlWV/wYSUFOVbGSMT+pBlJPwH1WGS/B8OBkPjx+b77c
Gmksb1LBILr7+MRTSw0GGXwDUPGrCeufSZLomw2oeL6Jvvry6XshgAMdHhDellmV236C5kgEX6Ih
moTuW3pTDfRo7FbNX0Bt2JChsLsKETKYvcczynkXdBjmXkpt0TGhlZByquoOZOHu/Pqnw/9V+Jd4
MGyRxDqYSMhFlSLAOKWFFPHK3u4qCFj2NYv3md5hKc3cinq1nWoH+TW6sgFoeH/XAN0rIl8Nd8BX
6XgEfWWWev9XVcFvN/D1XbA1yYx9I6zYZ5+3GPak0BCkqCtb8CG1QpHTQjvqtBkJuRY5NGbyzwuf
t70kEazJoPZeQKf5wvt/IPse3jirfUegTlBYuxfJnS+3yv0DjBWHMMVSS5L59N348c24EWqJohsI
QJ4+hTcasfLs7819S/eHmBq1aQqbC72Gzu5B76OTD5uY7saN3TjapgNqV35DSSCkMqHdxWMj2LL/
NpL1VlblnQZJ7mSdV6yXOPMmsGEbwYBoIkM1DnF1OjZbknVaOxgf9Qb4Raxlclx4F/H6yxUkkifL
BelwFjyt5YO2ZkOxbaq10nolPaiVGRwnxKO1BaacUkMlc7RJqgGHsNuCFEWboa0x2MUZVH2MPkE6
8Rx6Xl/t2t0182+vEB1B0SO3ueSOogXUcNsrl6jt5MehtkrM7VuwjBC2f3+tAKYRDDpZ0kIBGxiI
Bqpilx5i1II+doleMKZL3tCPsLx3KR6KYUyKw10iCL3GaK9g1fYPvKtEfnPaIthb/1uTEwolSjL9
Eo6YS2OBk/U8r4ZuS+JGAl1nO1syRyeoL0N1IgMd+dISI3G+jvnVXi9+IjyleFA70xzLPkqk6jdQ
gIR9jh7nF6BJyCrpgWeeY/bTWk+B0VN4iyGnfmEFiofeezYrHl4Z3OTQ5JCcUoKsSswkv3sge1c2
WDjVM3HIaEEmmdD7Dnd+gkCCuZEE6gOc2DyA5DWufry2SeEUTY4g+2FIaUUI2U9kSJJi1dP0q2Dk
2XgcSmsRppOUNiMxbpocy9Vcv7RkSgs9K2M7ufJBZhfTSBTXgrWBFanc9msf69zaQN5QxFnwHUFC
Chty40EoV1N7CGMg6q1VwFvLbu0dvQ/QQ40BvnW2wZfeOnzebiKIb8gKZdiaKQPDFdXB2sJko6c+
QCOLWt/SQ8ceRnIYrBF1KcPTDaoyufo20fgXtiGyQZM48IhgAQ6tkrB2aD3yuEOVLLpLEXRfWw+s
owwPwg7TvM6xXFr6paPaw+6KPGd+HpHZ6MUIwB2nRZz0aQlI5krhd9mlY3M7Z5ALFbS+lidLJb4/
7wrnOW1ibckfYeMoHN1CNlMewP9mHP/SUsY0d0qHl0KqrwUtmotRNTqs0aOnvZkNs2KKPUtkmGT4
+zs3WMVYlQHIsNaEfBUpHLeRjCXYoLM5yL+q4sMUgcz+DswY5zWRHD/YV5r29JpTIHHh21vHM733
BMCW/E136NNYAsfhzUQbYEPTgQ5b5TdF3xtj/F+K+44hYLGWlclq1G5GTReJEBbYnMfqmZVWteTA
yGRuGY5Gm4JihxWW57XaMrt7+AxWtVUSh7u7TNc9sFoU2YCsRt0ZCnxyP8GVAWxUsSJD8iwoZAT2
yDuyA+v0Zf4yV/eGAuKnSirKMgPQf569oCvYYdGaKkCT6bWYwyOeg5GAMJej+ZhiJJ2YmLbHJHJY
z8DbADVz9lM5UhYb6NFJoI/hC7NMmQk7nlHIHRu6bXoXkeLk/w/je4p3U1nssYh/21hovnZR8TO6
KBrFdTxDZBaK2NXkYr+AHvdIQZp533w1LDf3Z1sSpSoMEIIqIyHxZOFqs9FjSYM5iJ++zYU5xdt3
RIf+loHNaiQiwmB0ivmlbo6fhTtcFffUEn7Z3tcnIU2CISeY+mf/awowM7t1wfveT3OX1IPwfdE9
lCZc4aLuLPYxyw/P0NLIj8lZpYqNkhIWFmkzYamYcOQ1BV1ebKOlecfx8iUNyQKlgvfli7hzycul
jT2kWvKaADm4aitKIUAz14Lgv8/M/AtqcDIZj8knADYjp+ZSzvqw64GrF+55zzdFbAH6HW2cCVJb
5LipXqxa61rZSdmJK4qToKC2mWspaXZyR1/ECpRQnBAerHX0uH1ye0yGnIXjgX3528Lt72bcX4du
XZuWf5Vki0/vIR0MJpBjA+6xNa6XKvclFbrH0LxIqMYsCPbocXE7E/bS55cEQBEFbZZbJ1VZ3zMC
SBSjsErTUKvJ2KwZjCV+qQCpzbKIFUJsVD6u4TG9rNhItIddu4COQLExONdqiVm5sJtObLKBHOgZ
IMaUmCREa8jAUe0HeHuhQ4rd/wyRHpeURxRQ+4yO9M6+6Ba0loDBRlpQn2sRU046N6bLOvWgvJhq
CQ+3cLK/Yt4bAUHCZ/GZKyHOnzsvXU5eISfegiGcsLYX0OhrqnZJuhRe29ySzPVkECN12vcRPGPa
P7E6JSERI/9UR8Ya6aZVzy/riQ16OHKewf61L/ymcqc3I7ZifeUtdx/J6Fi2IV2wna15qpScqKCh
X2DQoy2e2WB+CbJXihkrzwYdaA0C0wzaDKBG/mwWdrohBSKHEsPzGrDLlnQvuh+7UmdzOZ9nIi9X
nD0lFQH4GkTxIgjXuz7sdixT5WU2VHZksfRDvdBSt6mgSkpQ/4yJOBsKRClXwRZEOnyE+RWkCYFP
Vecj4q83HOk9nCxktrS2Fwf6LXEMYmv9vcHVqHCZbsfdLW1SVx1TWlGz7xsWX6y0IzkF6U5ZS03L
o+tOJT2auJkBqVIx/mn6W4bZ/GCe4wt+6nacvc52tfc9xFCXrLiXt6pNUCC/CZ7uHYOS7gH0fmcF
3DNOvN1w49eGhG1rXMrD7sYPrmKiENjkKIlDEL9DE+IP/PwwJ+9olbz/9G4iLNqlbVjt7GdWZDhF
JdSnQBCcLVGT16apYelgGYiBJjE9aFaPPH6+nxhtwimpPjAJbyDk9mHEpcW3XqH58gL/Jk1Cx+8/
UEzTrh2g65pVpeYGqF6q3wps8S+Ze+/kGsQVvsJjYIqYEbNaZwl/fjWBlchguUnQxJV7NHfFEVLm
DQ2AaHqNRaLIWtISEiD7qmqyJ5Of44hEVDQV/s1PoYrixO96dMmjxuADBylfkv3VOfdlpraUwT5t
53dEHpXqus1+WwaKHD5McBUJXYHGUUP1MeqZUODABXbyL6/66mERNaXTzZ3jWsxiika48+l6cMv0
eUpL1IbJIFqIYUmQ18BurIsoYBZmsuiPn0Bu6Q+G4Gnu3iyFV40qCnZ5AMwfsycHtfqb9yEwhq5x
PqYqvVjDCw0hvnkk+k6nyXqbeb0v9oVp7qT5CIoSfbR2kMd/IRFxENMLq7G++9gdtF5eSUbGqcHs
XY/4vPRRggVYN861VkI/uWMzQkzZdziQvbAXZouLPvceF30n3x0reWfP+PJAotIegtFdi/1mgRqH
ASGOT1ui/iWECYRdoC0tvgeLNRm0Q+pqFMh1OCYtY2JWkU+YJzERrVfCaa7qFizp5YoPfhpOxDkB
e8SisIIkOhj4VskQc0vsurSYfWnEuc4RW77/f7bPGv8wnp2I1+oYPyPy3dqvtc6FeucXVjCJb3dW
SSxTwqeD5xQPkKU0niABUxYyjMkUFFDIR4wz3fQITOtywHDWIR2ha05lXPObxirPHyMV7HjmxtWL
WySG6xDqE5rCKL9VUHG7B8vSAvn157IrsOUaMLVd2d4A2sLTozsxP5cSJfnPgReZeTDwHIPY0V7n
QlvwEBoVfSHxNWDVsl8jbcy2LLRFE4YFRYWMi5IxOgRmJiI9aG4njllprNYTqtKqX+8fu1EZtFMO
EMj3FMLxVkAqUnX+nR/qGs72iUTxkd9cbMlRYRYtooLmY3FmK8V+cfyyqLSLgKOU/QhPy+pHBZHO
WpqHgWMYKUSB4zRm5Z9adKQwV3heUAYV4Cw6Jhz6QsUmiigwKtrXKUNukmryT+rtLUOc+dNqLgr1
McA+Ir9ceXsgiEbZvDPcUkbWJq+ZDs2PnJBWAxAkvS30FhznXBfrzJfFyJc0PREhU3dHdc8LnPBw
R1NBdWxInyk1VL6N1BHYb+G4XOg7jUVFBjmXoFIsHv3zmGhEdtPf0SGTlcWoXAV7aVmjJ++vxJhR
fmKpaF/SbAe44NSH0G+H5p2HZjFY05nDlEN62k1l1/N/vfsSPbYm8bxJ5+0/oEIFNQwhEVBgvLgb
s8oBaKo6UV5GgIvABiv2XofoYj3fG6zw8peBUqZF1x3W2BPkxnRLVhrIwlpOkXJ0SX5s8bnR3Izs
Tf5ZaUa/pUlcKdCZICijj+OrYzv2rIs0/cbxJrrNZlR8FiUYGZ3LZOrp/mjkxrCn9IygU68FBRPp
BMdhb4DIp4RqdHwv60INjVY7BsDd/Y5cpZcUEZbLuDRw5yNLNhvn0rIzCapFUdErOlAqsYxkmNAV
odlNhOacQOp+oBOv+MplKUn5F2cfFpBiSwyiJCbsRlF4ISzqu28na7cnplPEZKc4jtD1f/OM8V2D
bv3gnV0YhGwfX9z6Cnx4Eo7/+zAELxtjo1piaz5QQmhsu7J19Xn8ur+ibrzabaV/Jz4q0+DidhAJ
uCr7jN6ieV1GvUOAY1+CCqiP6yeXYcwVKbGvzSWaOuax+AvxlnSl10lC00nvZ32pDKOUxjVls55f
x4/hHZa3EU1Oh9ysEsST+mi1vsy9L0MUmzcAfpIJFfkKzamI4rpqq++KwL8H3g382CMAQczkd2ql
7fuOeVImtD152IkPrJcqP0tjP5EPkBE+yPBVZy7EU7vEIcGYo9h4GPBTESaMT5fQNSmTIIcsxkBv
41sVuVNhZiFWz06vt5KfLz/h5rxCEbqS04M9IEm+0ZXO0eXp+vs3vXqMM88YmaiV3BFrXfC6Mgzu
S0NGdUwRc+oLoPAV3/Z+hzcJEcJ9mC+d+bXd+9H3zhC++iNZmSQrl0/Mb5q+ODUfZsEH+sjh0Lcr
QJd7Kr4vTi7069H9CFNOgEe+5bNeLQJD6q8A5vARcgXevB1tOumh/O5sNTYYrPz0BosYuevD8+i1
afCO7YYK7A0ZGgT+oN7ke8YliXzV+6ycds6G4wqViqa2d1SOjut/fSBmx5ZvhulZsVS3xhykrxBb
LGt3btxGnT8k7yjNmoCfEcj2CA1G6NKrYR/6R61QdViqE6fbDSFZyEOT/5Ci8igIiMssYT5n9DRm
KSsCsrkY5lc3Y74AJpNrL3ce0CHAHHVT5amhLODjULkCLvi1UK55L3CICbIUe7f/fDm03LROggYp
mRl85FaD40YWacUtgZXRHB5VNGTYXQCsMRv+nDCXyda3kONvzqzqqXvYo64Mc7eNrUn6fVWYOGsQ
0XRxwZlle2nYvLvFcBHhN0lO2ka+6OZ8O7oC4JhP1BenF+PTh18WUZUNdJ6fkHZxXzZfSVtezGVc
Z0pppa/+Db+X0fwc22ZvrurpF+LwNRtv826k3+A6lGwIT0E89HLTZjRZAWe6iXLnW6aHfPy7aA8d
RJgQkDnH93f25Bh7KZHDzJrq5uc26YobVyAXEZsmEbiSEmZfDKnkTjGj02aw64QFTs56lonRCTqr
vhLpDOW5yeYyWDN/OkMwyr1aKixE/fbaS47LkJ9XC52ybW46MJrZ/HYqdJYkjg9A+G+9x1Pf2gYt
BEoyf8BVCIjFGgQC7SBjZ0+a/QQLe8VumCuYBz72lPDs392OEhhpDn1f4yUZpr7XqfVqThmgmRnn
ikZOu81VeBnCxK9GGIUZPY/Zr11XLEXXKTjn1HlMowyMRcqqShcW/4jrncVZW0pEDaNCENTewAFI
L2Rf5LLR9pv0PYgTmHuLmrc1ciZOTRCmRaefuiXURhfh4a/zKqgsewyx25xV3dzzrEzbPjtRI24r
TDpBZZHwRYgIz4z09SWmdASoeDJQnZjIN9MJOBcVKkjpfSmGAJOxYxP5HcZnyeAgEdmrVnp/aUpd
eDcVX+62IeAHKMD38cih4T8QbTF+yAl43V6Y2Q9bWWwaYryAtDZjMztXDlQY+Mo63mOGT8sakek0
b8sZtzBjMK/pLElETHyqm4cQpIoaZqfg4cFWg9+Tq0qMRmG0/vufbv2Q3xXM6R8ZnPW3d7WDJqvL
5AcXWdsEkUSmVDyHgXpDZ7hastgFnaVLu8b2ZQijMDBtY3TfYPdozJnELf5a4VeVSqQYm9sgrjKJ
Y7StMDIrQdM+42VHDwNiQ+ak+scvanMI69B6jwLqklD34ZHkIA7RBo7WBF1JYYma9rL3qWWoiGMW
I7mqfqE89aqXjXZQb8AQbviFFAYLH0hJ+BlwG6l7P9faRl8vBrUPUYPrOB0ANmztFzC+U5YXue9B
hUdFsmzIinXWNEH8Fx7hzdeGdfrZtLOstdQByYpJGfXqSXGMWYuQ2JrqWGOcNj5LAvIJ9ePvayen
9HJPnxjaRtaQ+kSGNiZwXeSazB0hGWXXBpF7H9YzWaD/qQtg7GlwTMzvj49yeRyfqg8go2Xl59C/
fahY3JKpNMTSwhwkNyyFI68u943ggJY8gA/UI882deuFdfAurSxMdqepnncr6jvi6B+weqcuJED1
j4l5BI3s8LZ3TdUvdz02r4vdfht7wxX4GXc0yc7Gr0JoQIxkUSXIP93GhcHrmCiZG4mxBGB6sa16
uY2A7an1HLQ7ZiLlSgy8vRTfxodzmq3SV4z0DTKjKjdZAVLOwwzPrwBX1SNY7oki1vkTL1V8ObkZ
+8melDMzRp2b1upObD/HdfM5qbsoYxez9l/zfzQIMQMsskJVAvhZjBdIRMvR/KqQrQtvSCw0+c2x
JAbIfPPVb2EIbBqEYzR8X3BAVt8n5VMlIfMiBv+epXMmyviNMMGBMH3QWQSgwVQfuC2Z1xAaXEEL
XZfeyZjZ6uAa0tBHuo3bKH+H/sEWi/pwxnKdjw60Hy27oFVo0nyswmwWobs6TL4gnFpPNn3mUSrz
zoscZavy2tfHTXWVTtGHSEgz8IJOeg7yVq3sYoordnSFGWWtwMciK6lRaMJrNoZbvCMntxe5C2vA
mtG1TWg5iIjDEjbi1XPxUmooxo3lnQ2ej5UaDNRPHwD/kVpJyhSReXcZWIbmrYKT2Y93abcXa9s5
a9X9qO2sBsCC7QtTugODXNYaNLn7WUuJJUdPx/0rJHOSH+87W2LS0tImhnLNXwsZmmikG0xS4OVl
RwEub/IO80SxX6H+5e8m6Bp2Hp0Pfy0mEI3ZEF6PFkY+Ev4zwk1vs+Krhu02YKOF7DsOGMWA/iTz
zwa3KwI5CTvZoOVNJUMPO4KZLky348oD5I5Orjt7DuiEsuu0d3IojIG3+rp55nCmYNfTKctTBQ27
ioaNdi9cxPcu+lNVTllwskhDzH9GtTtG+fw41bW85aaLpb0Oe/gn8CXvOnsCtPXh8hMs+5/U1XbR
Ik/NtSfaCKyxAClPR2Lkeq5yP1E9eGaYFFCzZ0icnnXNbgMZFwlu1i30CMpIq2Onv1cq//hCFZ7+
jUfZEryHG75Oc3GDMvrZORWEV2WR351chOu+9eAL5WLrCjpIDorrsbJQ8zU1xCpPJxAugfuKgLsm
0YoJm5IvniPE8FeHooYVxxz0FMjAEvppP2HuvmKxi4xFlIgt62kYv6n9gET21TizkS6BnnMLJY+7
lf/t2G4MPDs3nqWT6I/2aDF4fyycP7Z0pBATStnFKsEiQES4ESF/gBMBpjRtBAP3XQbxdo4YEE6L
3xs9sSr/pZGPeg1iJFcmc8ya01OGdZVnYAMrBOXnjJtLNfO5qx6fhdA5PRBDxpDdf8QRXuU3WqHo
wt17AGLjQRYtDKKLre3AfE0T+hvUBPJsEHHUXh0S4oPX57vw+LdSGiIdzyKcosbJzNSF8rFYGLFG
omxJtZwfibpc3/mpj45G/yYprMCEb0sszguZTpiy+BSk7SxIy6iWsKEiy0dm4Z4gUdUgUCGw5KeQ
x4VSFsObuMgE6YqQeXqeO6a6s9xhbRBsyekPA3fDvHLIJtGbRTPfTAZXHjARlMXs5suqN83RaYiO
dIzrlubaGE5ycvCJYF8FUZGiDjTohwmt+ZT1XODEf1pKuYAgQjI7sCPD2a43j0BXyfKjBQyeCBT8
LJHsRinACM2bkGGL6aRdEtfe3v3T0XBwfzkRCcSro20vXqO0OwkM3nS9kNdMP4/UvUt35F56pOwz
HfYRVatvuocpHco7YAdP63RjwYRS2QTIqVTiU3aoWRCD9YZQ3wlUrjQlHQAZaV3Gs4DY6jFAWaxG
qlPaINiS6GBGIVxbQK/JKO+2GaQNVypwVToX+/xvv/XYWp/6a+BtnBe17XRet/okb1jYYdehkqhS
cGKHHodd4rI9RC6+mg+Kz+89+AXJGIO2xQa5H19qSZuXZT2Oppn4BJhmn9I/wdQ1UuXEX3OeGWZT
Nk4kxcQJaFbhs6MKDJsKJpjMF27y8yJzN6Sly5uj4PJLeMQ7VHjwupq26Zmy3HdtB3+Wqbco/NcL
uOi0LQY2QxmvY3EhFaRxJLLUL+ty7/MduDLjuyoGBDRRtg9x6nYtsRQjmlaWJh8Gyx1I+Fsbzcn1
SNsXrI5vvrovDm2JjQDtEaNeMm7eX6AuotARCnrIIkyfXrO/evFyVX9kTpNGGgo775f+VbNAjU/R
BUCNj6QcSC/inna2r44X6Bs/l+0YwnuyWeC8zr1f2tJoJwTjFlbVo2QO7YbKzO1xfgj9crfeBbRC
ctQhCQSiGsdnNqrjDuRgGqTLIvncvxYRXcroEwyfBiYpZ/4ROy6wsvr8fJSUYz8QwjIG8xb4B7cc
jxkLPESQdmiyxw7vMadR2wKG+9lnuPuLUg4P9qB3fTyczttR9ZKMtjPsFFGM5tNHry/wXGTJ5WZo
aZnblbRUEwjQR3HheGogSCg2IwWE1LktjCGN3KTAlkKby+88NQbfjsDZKaloHDvo8bxw6Ba/8CbU
adRu19Kj1XxZZElFzLSnXSbvjStvV0jdKSOBbLR5Mdv4xByf4E+vihwnedA76XjOZRbXjkfv1jXP
ckCGxXuTOAYy8TAfgsyyC5jJt3POrTcXx9VjoJYQhur3mn60EGVKM3ban22EF96lU4jn5TsnRRA6
2WsEl4xUdW9enEtYRNd0hYQ7xRLaDuE4l3wWr3kkYMN0nH68WwhL5+ejoxk8o07NLUe6uZ5m2uQt
wYb0nUCNrOS4pXN4zG02jJcoXRZhtzdsGgnvlTCoofv6INOmnRvSpHGypgytlWbuCsDQIqpArTsa
RKVsH4Y/35l4eo6/X4UnHVgEeLujw02RbXr+EbZIPTRvKedsK17plRlKIq+7H4GIkYWAPha/1V9A
7J4Jvv3k8FU5tMja8mg5yr0MQoGgg71kVQUtkn4rkaZb73e66dzpuL6sFiH45FlwydlmoojE9GeR
TMBhl9iRV6oUAiGC0R+nzbHO2Qf1g9ynZSC26ot+p8c7q+SQeZKiKsU71k0a7fiPfg7zkO4hmW5r
33irFdef9pz8/dPvIx81dDomzbs7rjC86aYKCeCp9oEA92wYBWLTvXPIjosrtw0YwICV33t2QIZ6
s8A3eTwYanMv6jOreozp6Mb72hdd9uibKiC4BFXYqjNRaRImq8QuNdp391F9MQuKA2gGiDN5NGUl
tXFdrDFD/ZWZIC8m+S7dslDJJm9vOMowuxF8nvAx0hYkh+b/V+QhPgsFpwFewvi5TcxzF/svFdWc
w137Fg1JAUGwTbJJ778KmAt1AERQB1REy3vtkEES5sUUX44ENN3Y1EvdV0+OC6cqGH9SRWwROPVJ
wu1pw8hZZLz1+FRZ90qtCupjpFejjZxDH2X5M704ru2oNWwBGnQjFpKV9bDeyJM76GXpRq17mqIn
Zdgdb3rK5nG5bZNbyXxeYA/vcI7HEkRqyQezkeX3srABZgxRRs1oNLWpPdRNOhLHqSCaToWOdLlp
Z9R3qoiT7aQhhbFWGybuiZEEDr72VVqgdvVPdc0ZveoTRdKbHLRziyjUveL6fdVSR4IOzXLKxdA3
xVIOWpLpBObHCbEriBfxt+neNydvFREiaLSpIwmG/M7VCzt8H9CbUvK8snDhmJLaRIKl2cYYLAU7
ePCDycdnExJ2zX2k370FuhGM4I937W/H2fomlvuuH6rFm79Cd4OCEuK0c2iSeqOk7pdeaHbL85CU
2v+C4Wt9rpUQoLRVzJIeSoErD1Q/lOhk24h1SdITf1FaeXEWQ6bnNQ8+yfmDzNutULIkGX6NXP3+
L+6wMXMZFPEuvNOZ/qHimlH7H/8eOfeyjVF2nhmb4pyzoLxGNJ93YkgG9bAbQbKF9IZktSdBT3ii
2l8Sr3pVr8sv/I2qCOlJD62JJFoPt8Su6M1xItysmktdSuvj9UnqcjOPhMv4mUG7AATP9LTIawiJ
etrb9ZpSuO/UkJ23iUkrmKG4525Oin2pYp+bS+4392Z/E/KVeRzZbwLfQz4JX7wLVvmx+VmZT0AB
ZcmB3+vdKr/JkNkR0xDV4eDVfB1O5pIABRdZWMpd2ip0XqRU6vh9oO3LkoPP+4VOQod99bWdKHqn
HXO0GsH1jUgMNZMgtsWEM6G8EPO5Lzx/e8zFGXxDd8P10L50Nzbm2QfQDwFJb/G0JmDdWSt5EwA8
WD4+omKHy4MrME7tu56m9VZwKPISDClnTtHN7w3DkNepJz6GFznBjV+XpTfBJQAhcwRluVJadEmO
EMT5U7kQQYMk4QRMPnSIIEGeYay3MKResaXvRJZNqLna4OozFUvsBbZzpDPS75fMAEkSjb38/uO0
ok5YBEOGti0Jur1LrShlfTFZfy4liP3VOG4AVyAwhaI/2ksbExlMDWr7tav4X4tlsJfkJvKIqU0w
0gFWCxwvvV3qL87ZTPYVWoUcetFIJICttNqmw57enGw0SQPs4TwvEPaChcL5GrJsAafArArI2Ux6
2gS1OCShiR3R50N1lun1FDPfFckQfIZGCXaI6M8ZnLr2Ge9VZRznGbBpkbgTyNyh9yLfQVD8ZfJb
KvryfrHrOMBKoHNFE+JwuXHYlPdA2heyG9dxq+ubW3fI6QDLhQYuah5hbf4t0Zw4s1hk1Gmq1357
XXxLaQiH7qAqflx6fBGXVNGpfABc4BEmjAlyS4ZTq3PaMw+95vLEN0HM6/vA+f6i9LxJvFHyIJtm
SZ3eyLntbX2IM6Vq5RWcej0bj7F08cQwC5L+xR33WOVVa245g+uWRGnthPTKSPNhadPqGTaGXfPM
35liceQD0VCQM6tDpFeCjI14iVcnb3ekrj7OG81iZoX8fx4RA5iK1bXTHiZ57ests7/UqNUnkQaB
w4CzEpc7KY/DjANsDv6WfDEkTfWImtXGW0BBk80XPRpPHXTS10kZAE0qi40BqxbJ8cznH0pKHyLU
S02qsrxY+63VkUqgL0BS3cFWsS/H4MyyPEcO4IeZPBp4MuRjXNZH99NyM+R6weYSPlBDkWeq4spk
HnD4OlYzBy71JmUBWnsBr/GsnO7ZGDK4stdq57jsM7gw3gWXksW1kKzN9ZPHJxNXg4qb6CvjFAM2
eFh29WFpzI9cmbiBW4oybihZ7XpbH14bdzyd/kixouZZopN9gsB8d4U7HIAA3r2lHfmmUXgfbmMr
SSSdW+RO5tQp+rB0fidsueHbePhpUQZnBz4zd08kyYi+x6fgsRltckXMP0nk+H77WWbZZzbfHVQ8
JLtzwrMsmq5oHFDlkVAmIX5zDuqxHRlEvwptt2QuVXOoxJKkdJdzebmvPD92fFhgSrXqKpq5yBpD
9px4rTGJuqbtmh8xQg27bE0Rt9usLbHSHcK+zXBCxc/OWzZOr1LdqPSTPOFPaRkkzZHvcGUSw2tx
CnlrtlEO3WLoJjouGwmwj0P/Gmm7fYsL+XyF7wqBBG2J5iw6Kd64PupltfknZkE5JsvqiPmC0ByK
c3fxqcnCqsJ68e+Vp+ribfDDHCtE4WmhFm1jIFsjEok7G5JNvN6e1QdApv/YiWSoEpqw4+P3jjZH
67yNQGnetffGEteE15i1Is0qSqqpCDlDoZNptZZcnbhkHDFdf8E1r160/DoUpJLobw6pIflvRG0x
ERSb6CabdJTtMSlMD7moV/LrzKS6EbNzIQX1wH7FOF8viDb9AM1FVEy0n/N6AY3hIRDIAFhFZi/o
/kr8U72czDJ1rTANKjC9B3EBPeciOERwrGyAOY+Av4TlVN2a2xNnuUVOl7G/TDehYgB+bClM1EXh
Hi6t1J3H5dkn/nMr88MxO9vcKZK116+0s9UrV/IfLycwDB4aWYKhdCfMBRHNXo9/R4dGqpiwVHLs
8Mm4N17a7Ne0SRbpMEGaKFdTQUWEXJn0/QrlCH9aW5XY/EnwOqrwn49sGiK6WxxEoXxpsyoy2P11
z9gLHZBsAQ0tf5APlRzfw4fF6nWYIgEs4NHPPQm0DfLIXrxezwj15vwWGNEMDYQ/CD17b73mgLWR
NyYzPjwNAp9LwtidyYkg80bJ8WdFRpyflbzYbEp5pl1CV2SKtpHQ+gnZ2fSTDShOiAzBJo+PFHyv
pY7JPug5nywXS4yeh6Wqpxl8ZLEIMWE+pf1q+D1AiYWX1A1JUiIFpFMOJqY6/p56f9CbmAuEfEbx
5wEc2HmEec2t0MYSaPtErX/KqrhG57h1iqImqDoh2aSh2ipwn+jU1JtiIZg4jD9u4pU35ib24739
7oTA5Nh5h+sEL8M6QLHlC/7XHsaoj36slkW6Xy/dc0/bDY5agR/Joi5SCyLvxS9nlq4hFj+X25n6
MDenM2Tc77FiwzklWVsQVIZ53RGg+vvTXjBHgONrquZuJ0wyMd0RYclXfsoySH2/Vv2n++MvGvAF
+1/q+kv5Uu4kPnhPCMv56TIuPn8EpiN+1ReNkOkpYvMkMmFOnS+EqsIj8PjU04UUCbwtWkHx9nEP
qhtHS5bvK/Ap6GURG/5EfotQvUOPB3hwnsKRL4iuTyJtARKTXN9IA0pyp3+xI2xu0faFxJysOyqQ
VlNcWkBvskPCYe7mQnb0w24gUr/TBNYzSB21VMiWwNokrswFg0EZ/ykQ0t9X2pqxk0/+qvh796yX
5+t+pGZCvm7Y72FTSVVx6KTZBDekLhFBkU7gjBCBFARvOBRTNRTsW8WF/0V4Pzib01LmSlRavsg2
3ihpEGHN9B0TkUhuIla+hA3jLfuspH4dqNSS+8VaHi/V/vDxF36DE5gcFfAZElaWtiPzSZ0tHaqt
YgO6bc2X17EMshfljCsYiJOgtfkNN963Q7QN2InJgRpypkqoCqK0LZi95omIC15q/cKDMcFbHZ+d
U7qnLu0xw8ymOBWTiF93NPyNUh+PSpq9zrwzaLmGc5oIBcyORU3eZe59K9V8XwUnR4h62j9HalUY
+m2k3ThzCI0r7yzDGTKvxNpYK+Oqngx7QIhBwi/nEYNrXNvPL36j6Dwivx7YJwraaEJUlLDmnUDX
Ak3/jZ4tnOcV4KJ6K/Glh+amSPDFqUb7q8Zqo4euxvvC9KVpPZa+v90Yip5xksFmLH/rpUbIdswg
Ehv23uyMc+o6q482gwmMuVD7VoelDimLzRbdpKwuSHYJjXV1kzWp0pNSMprT2IDUfJVanqIo2YG0
xu3RpV3pdOgLLM6WyxE+60iUDfVWDVHqxp0lCEzJ8Yym9JKgXsUCpUNEowtC4utdsLh6bGqrmowB
La+FfJF1ybiDMaL3Xw1HW/ojmAFDZ359lO6oymIF2bguNNzPcGjmJKKLfU8uImXVAtu3A8XYIf7S
qiubmSCWA1xvpZryl4uPfdjgw8WStYCr8q3y+QU9o/abqB+0urLCIyooEkCE+JwO3jCvxpIYV67j
xvTsmc1CnqV2woawxkURXcelIgR2exgrB1CkxEc+UQCo8Se9G+DKLp5ZmtUxI8gQnEr9gH8+dD0P
8yyCqMTiDMwNBG/BvHd/7Q878T7zxCySv4EXkFIP5fWCc1Wupknl7Ev4+akVNT9p91YGCc5vHV4O
wGYGg6OTnHVpwTRhhzaJW+3coGhMKNp7ysE3EuXzjGEzCKCATNzM2X99LqzmAgA0DZvMy/o96L2J
owEWThI/B+sDNY6q9t2E3y/HTwiU0+2epG7cROFuf1eL/EInoieVLxPjgs6+7Q/9ew8dk+qf2mcU
7/CkEVbch5KkI8fQIdPkDAR25ZVyc0K8EKJ3q7KxEefWd1lclJciFcaNYoRhixUakSzAxs/X2iri
4Wc1DTpUb1981+Z0dh+NZTeb8wXyrxvOTNQ64BenMDhocCfOQOr73wV+O1OAUOK0cpV2SZKlp0Gc
QJobeYaNJTJILtACGTZYNeX/DfrnXavu/0KrDrVgQKqdotCnngDz6s8OW4L3oLrzo6b0atWeq27v
+MnkFjytYHI3vkazm2WFZ5iQEwdcRGDuuxvHYmlQN7oqJMLr1V8dfXISlnrFpd36uo8nuoNvPddp
jU94nJfU2PuSp/Z4tkd6k1MMsttGj3ummWpYITc5S18E0Tu9YBzqmhFQxMqrH9XbPJo0q87rJ/pZ
E0k3H8C5H8QTYp+acJHu5jDRmpJ13yb8kjHtrbx7hmuGLh3/VUEJwAQQ9xTJakZY58pN6dpWW9Er
FJ+/QN50tp63f5Qb8W3AQWPvdaB74FpLYKHPOps5qkuXy2rdY5+jixIhqolHtewJTraU5QSxLu7A
d66/c5y9iOWukqqV29IvyV5KckJBwPFMYf6AuOcOUINS1uN5il7MDTlw9c0LfU2UkV9el3N40Bx5
R4D2UWvsUJjasl97/dxDVgB20WkVyPtO8f+b4oITz/QHwpwH1AZzTag/+vtZom/TkNzanmidmzOZ
n6ShLuZ/jBEufYyy1hNuTN2h49fUFzpEB3qGoNxBFRjY6POotSEO1bwduk6XJo+CsMmnPnXFcBfC
DJwbj/FMFGS+h98vQeVlAUvBH3e3jNu8cAWaqMiZ6Em7+KJP2qjdzM0v5ALVMla9u51Kqf9ReE1S
n0AjpvMC8jtO/k99229FhHtUTZxxh/ngGYt86q/OmpoEmLEq00b6ZTTOK3uBvyZLtXFTXG8jY/GB
vSFxALktV1d6R5edAP5PNF9TNJUhiwkFVnIUoKWq9J+uOkz9LP+3eaiJR7JrtmvVV6RND9jEq2FL
ftfHTcKi4Okyq5Hk4B8q2esuH+ibyiBfZD6wTXgCQYqcyKyTDkr7q+IFVfpW4ExupRLfVNMCtOTx
aIz2QfwPrrrtjbX/NfRy//cGhZQTjEIJkPXhFupvjHNU4gNtbpnV9Vg8V9vPCGuzgrzTUonCuy5s
ZFe4l+Xx4NFko5YlP3blOvJ2G+UdC9sNs8NvW4BwfET+a1KFzx+BSmQmxA75u2GNloy8an6qUPBQ
TDURVuhgR0CqRcqMnH1OmJZ1htaV5J0ush8qxPYsEShhh7r+oSTOy0F7AAOPvYpFU2naOmKgV57z
gUgh767iKWzJ4Kpk0HwtIcjQFTv3n/u/CyFLVxkGkZMNG4Ifk3C1NptlwuuPUOXF2K0zkNETN1Nd
6HmgT7K6De3Q4/lc/uTzKVOxZU5NJ4MmW6T9GPZskb9Bq4eaj0d66rI2B8eIs3Eefc/q4LvRh+S5
Rgo6PX5qY/t8gY8ySwyIKaasfkaqi21NyG2SIqKFg0ndrmOKB5fHbWN90zqS4h6SYzVFUbqS6DU8
V7FX45pTMndYbaBsezRQXwWSBSiQisQPHXe60MV4im9oAzZ0oNuz2m+BaCxbIMUvSUNGfZmb9mio
HvkYo0rkjCcQ4JyOHNgy8C+rmIj+hDWtVSvDIkQCiGn+HJK7jNyWryBvsxO1KDuHXjkZ5UvwsMFj
VP6m53sWlHPPEQkMdJf9Z17nJeQ5pXU6O/PmKnwUsoGXwXYa7aMXYAW1RMOD0yR5zucP9pi63mfG
XOft/H+/THtfoNl2gKcrfqdNGP+zt1Y2Y2HxZzBQ362CSe2Br0Mbf4+Eqg0a9dFiGTa/wSgnwBdk
KhjGck5W4IG87dEXVKNpUHZ2KRu6RqATgQGY6ZfjMtj+v33u7yi7bS0lQzmhenPs2Eyo4ZtXFT3o
1L699TP4gKEN7jbY2XRVmd0ZBrQ4K9oS8qxUV8FJRlh/4+fzBxddi1aHiJpKi4Kb/nSzLkrT44ST
PPMRhmxJC+HJQ9lGz2lLE7Vp72urD7o7e874jCzIYoS17m29QInjzlW+rz+VTZB5aRED/O+5Iter
mhyvTS9SKuFj29eV6TO4nW/qKy6dPLgJMhkwWGyJUqPYXIey1puWTCPu4dr+wMnV24vfTmWs6qvD
u/hmjzx0VbXLuQjfHkC0vBjj98Gg3AuzA3ICdcahCCq5fB3x1bXvRG4yuakMXLVvpt7BfWMkau9C
ioMy+xqj7ekx5VSyGjyKlZ0s8qqonXMxrV5CWHA5H/Vt0108zCqk/9ptraql+fZ4vLQXq6QwjR6Q
PHTsx6hIYNu1jloCWHNjNGzo3X8aVfMFpJZgEI/ft8rcBRz5Bmmuhs7ZB/7pPEVA8uBd68UWoaUd
1FNvoHVLdDcWoLo1Wto/4DpRIyePlVOEoFLnJI+nVfpFsOQF9ayzyRu0f1+USGQDZMmYFjJQOdVV
czlpXlPRUupdbA3O4kE/59YkFQ1yVyMpkvNT2J8yMtR5PhKoDLCQcq9NJbZFR2uqstxbZdeeACQV
Jngp5D+COpuqq+/L5gDhnZ8m9ibaMkJFJddiSPgBka66+yVPemcZcqlQw30m5acK99mmtjGDGwnv
kMxfEFiX+AunDh2heJNmG1Uj/CL4ooHXSslkVktS09VeG81x7byfzvBT5fmPGQegWtN70b8RkmFN
V/e4wtEdin+MIGKJyELcYMtRjMsx5S6gDAvjGaapsC0YPdbjkKvH1vWaA8yySJybwy2EgdRrRRTM
p48TxqYDcvxbPltdBa7Y3wrm/UQKao64qiEq+HPZOoAOtyOBXmYGbkIa91Ef7dm2VJWsz+BL33/l
s8TWgjI1WYk2jLB9CQIGE3Exu2dzvsil0u4KnsoIL1AAHxNrSpDhyfr7EJnY5HGVQyxhVh642+h8
Xk4rK4N4gkNliv89DzSeF0OPEKPFxt5/Il8qFEawK8CZkCjfEzL8kUAprbJ8uj5zrivWTtmFBt0B
AaAa6ONNSwsNCFiKbgu1OvrrMEoH/XlYwiHsYUA6HD0IXPQRyZKdKjjI1y6ImRqM/Vfv+YEf7WnK
3KaAE/0y6C4zCDemZClWqKx+1j0D4uZj5pWRkMgnl9ZczZ7V/Q74ODerbvqguxJeZgaeit8Egog6
N5RakqDQW/77JycfSNkainKetgP/D40UNw57Ak38M98DDNrGVFVelT7d0xwKU46pcb6bBwCcyjbH
qNUePnCTg5nEDQI/F1Ukcjep7Rpl4EWto7dRuKoTTzMK7gmgiWhFFoqynZINNAFB1qR63hXJga21
cQYRE6whRM3rPCIqRcTUojq4kUVLxChOe724GfdD49BId4+9AhuHPdGNoekq7nJD5poBt1LQzq7y
QeB4Z9uAYDwJyMbnadd7pmNa8z4rQAXt9gHADzY3hRMuFKBwTnPxMUvCFCongv/xlwli5T4bXneH
yuthV8qxMC5TpIrbWhIhz5EpmkT/IgJgbA6mMP0gmkjqDwjr7hXGq7RpjUWdXkRQGzGInwhGy5/h
TRMIx8TXd6yyWvnWcJkLLkk1O2vB9l6KldGwKobaiQKdEezdSub8D4jdufO1DatlmEIv8YteUFVL
5OSr3SlK6VlgVme0nDdbxswK9TbvVVC67ACv5trv3IJfyMuu2lkoqjTtyUeMaJdkb0o0cKswUd/Y
qCOIbwVPzC3R8mUPN3XHBfma5Gp8mJf4bJDQY8lIB8IpBfcq1zbC1BU2+v5MSQ6v8/GEJ9iv3NMg
xxI/WcNTsjDT5P8ACJ0MSpebe3c1664D48qXmJ6XHOmhf1nOIQbD+YiPRQDzKGOY4CX4bjRcsrni
Moi/qHs0sOwfHPJ9zVR1DnNTUdiq03D7X5x9TV0JI0JAmvNops013+mD+9+cqA4uNF7R+XhW8mEy
pKuPRCuQ1UAbDSqTFU2X3/OS6aVfaoimP6xjsjvk5+6TGyHKEs3G/a+I2mVN/uhn+xiSA57DifOH
ZpQdE+DQwHYBhe7ykUTOqmCqgB26GZjcaQDflhKqdlYju8TdG0HVAeVKVkb+c4t5WMRiDb98bZPQ
niKTsNjo5m12oCWi9ZjnfSgUxeGYdL2A0JnFfGqUbHEYrEOs/H9qBuqaaRTtQ6rAZr73gd9elChg
qAnHZkpZMXNfEl7wdTcvB041FkbtqA73vSvfVMMPpobmkJNusIHfYw0jaK+KRd18F2XvMcnbCJMI
1oOqydKbJ3Xz39WV7xREX395Kl/TrG8d++7EOY1Zo4ro7/UtB6VZjkj90FBmFkM9blcIx9OoxKGi
YffZr+LSFnN2VDTaXNyB98YfX9YcBGa6/EwE+eBEd+OYxehWbLGtzcnbs2Ws5SD8CMDnMafRkZ19
Fg2mCp3r2VLkbQ+x5/iU/WPRYSLhXQmKIg5YAJz+n9jGj9161WwPR0RDrBbc7lN6tf+g2+bvyiqA
TTCDYNeUryUjrpuLeU+Dp28JdwqfKXEwkkb5EvkIyQguJbXc2ORO2VsgwPs0jI6cU3F6Qbm5GOZW
puVi4uKBV0OQkBzMJmUrjrVz7j+86oBFk/eQfDZhOZFN3N0WSYyWtyTIGrD4p3yubbr2Zjn69CEP
ygNdRAjlJNwyxPbAuc6mzsuqrddoDTdiSUDDBmfLCc4K/JeGVMwFCmKpzfID+jJNt9JFEsUugiA0
tvbQQ7hdVMjun8gz+K/0jbyf9svwkLw62F4dLgwoz4gf7KGPFMzXJB7CojzkgzLRZTEwwyb80vX+
ZHELa4dqXI77jjyk5khQIv8fq2wVwg7vR2CFmZwR3QotNmwr3SwLQBRxSFKP3EBMvAuJV7p9ZdLj
Z+HcEnSeuiXWpXyaSh6/D/lkB3KkGjBlE9mJhWrjohEmoievWVuwTcDKzcRmLvPlHexDJErSLSbY
HOtYJD77IBOWJ28KSE5nkOHKIK4ES2vsxXUFMLrP4LSaRsdIyvemswkS4SbLjCNRgESCcjAJKwMh
NTo46PT3cl52iumJcupDg+w2+MbT1k2Dr9Yj+vKILXWAQ3aY/30b/8Kbu29FrnSoHcIGRjGWeX8Y
V5y0gh6b+16ZEl81Jn7SCey8xPYzfYVAKwpSTnXXukHbMXmELYz2S5vt7EJAIfP5qcf0KVdOqxZ1
FSQPvh0QBKllf1AizAaxMcu7HBYbhgFf5QZ8pmpVnzGtuN0+OdTxSyAXQVdyMur350mIO8RT1Khd
C51uL9jXuQwOZgHpqovVPvA/6fg9WfmYCdb1vgYDbknWQ/b6YYY5f9NQHMvJYsL5bT8eudPOsWnk
VNUrA+LmHk/Gk5XAvwdhcUBUX2Hls3PktVG8WnlH2hSgw6bquBGR3wJfDXm/GMn32OrJNqtcr72t
JoYawMY6fR+vpNyM9aRMoA0sGz7+o/NpZoDN23jLCraEI2fU27oYgj5a88AVziYvKrDYF5TujwpI
np9UDYbipDpTTN0Lzo5GCfBKKZukCwNpxqMYvCVbPOCY9SLyLFWoE/zbsG6y/6Jb1CRDd9x221wl
pNcqSVaCvBFcH1kAVI+a59vQ0mPSlFJ5hrurBFX1nklTD79+PyWAyBiS3Lzf5Bvzej7DdZA4rclT
J5aOB4yXZE20mcTKeMh5q6hYkOPmEqAjilqTphoqPUjOvPWo25LVjFStgzCx2PT+aJPLYkih7BTb
yZ75UzhkRjUo4DAiIuVRIPTT+t3upL5LrtWEyFCLkSbiA113A8AJXN8p7eL9nyJedut+8iFiMwi/
fIQBpfmvC3yxxx1H/AeDIhHOuZPb5F0UDjgEA2CobieodElYiJFrtuqWuLxjmlHIgFHyK/Fhe3gO
ChHPTO9HpGHDwBWmMXnVKi44OFAf9TU2OftyWRc08hWXEHO5TA5f/s2/e6fVjWg9R3zId1ZBiNCj
YL/+Oy3RX0bDhNxWeRM87A1M+JF+lzvkR5EnzHtM+cM4YYyR4sDtoW/BH6+/4ihuK5AlRgsqDVUe
pNqY4bhIcaSNRPyPROLHdD9/6Djmu/F1BVqz75NJhnBpKeKSJafhRcdG9xHQVBZ7NXjHGNq1SGo+
jn/tL3vyYCr5fnhZh8U5tlm/vLlWgF3qF6TuvIX1dmkq5o+9jKVkVrHNYOL8P5l8dGl/iEaoZeo9
KiA9wF52LePQW24uNv+qdKXN05EqAzLgVS/IZYCoQUCal+H+pFl1r0obNd53aLm1/P+J/rlLDkDy
+2R7BB4BqMnJnQHziwv9ofmMBhAYnlpo2VP+yP71PJbLF46ohPnxmfJXd4AjUGTBeSXghGpHftiN
alsnmwcUcgy2b7JbtG0XI7K3TFw6+cjGd5CzZvKC4k1oQITqCgC0J3/cjhgMBh3lHAaoQIFJQ5S9
fXxBvKeqyFqbLNfFbN9NVE4MoHR/cGx02SCsBsiJ6sjkOd7nBPTX3QnzNEd3nLKERz5dwGPgwMhQ
kU/9CN/+hzSwfrvadHh9cLsA9NiZmgZXwIO+HKFqh+xGGmxAVM/kYk80NQ71Re6/6yrHT1dlSEtC
DTRRX2cpQh0Aa/YGv5EChkEXEysLGUYdNcnuk5xhHIYf7RXz9i3wBH/PjsXuY5i7zb1ozyEsJDc/
rmUwjRI5F6+YwgChbWuPS6+aF16DzBxzlcITwhhMzWA5XwhOpBKNG6L3vcO6hdzaRMZRTKiNEpCO
bQ6NX6nvVq8TsDg3zF+UHBjN/MBOx+ZE/W+OtKjqbAFw5r//c5CBZBd3agnM2c3RFJyIHpG/DQ3Q
5RLIqzoqYccCt/DFCqiLtAHYBCkaIihKkuuddCSRwmUS+cSwvUPVRtrpC2uO7akSAtX/XKdduRUC
GsyklHrnNjAn/lZ1LbD2/VguiAEsYrHXlIBdXa2GoaJmVcvoW96II8ZLk09IZyzGYh5bXybnx5P3
zE2LpcYXk+gN88Y9X4KzO9RkTKSzoanBcVOT2jfAov7tZEId+o+XPrRIAI+SQG8RpLvjql0pTeYe
XAAH5GyxOjzSKsvXte+b8EFabTX6dYiPlPzmoIPvthoFgU+yauG/Wwn3bWpsth/1UfcnnR3tASpM
gCxw/7qWOYYbP4XmJk3Z0AKV1ZbKeBWWtWDDytJjFzS5jOctnlY2CvJiNSncviJA0MTs02TBxzhK
FeoCXvWgx2TpSzWwWJ95XOarasXaLYL3wNEX0mqc6ASNicJss912uXllyPm/mBdMH6pXL4q6qSZ0
D1jkFeE5xphjhXWnCkdjZ/3lRKzKi7Ztzki/QFp2ylMlKrOZGpOrLap5l0v9SBxF8nJBT7R8hPNh
iA7JyFwWplO4H4rHkXYQLuibZoYP+x5LvqXzawKgmRw9149ktDeAEjkuUFgBzMzq2mMobJe17AF9
nfe2fA4YRt5cxtc9rhFrT9T5kq0BvIB7yHhzOcwnxwZ2LCYrTa2hjipm4y5RFJCfwWra2iewm4Rp
86G/p5vqRpWifvrwdV7FOE81jFfoGqphiPrdvi6Dy1TcggfMoxeKME+H5z8UJobwv9deKQmzt64P
NclrmylxUUQJjlJQKJp5WcNC1n9Nd+TGUdd6iyMAHa7XlEGJe+7ywq0MULnoYVwVcw4fjyPUwMK7
MclQbqPhGFovSRg3qfbM8Lv6AQrXs+Z4IKm09H3/arD6hWxTcRPrDFersaySnZVH+D2TBncnKM3F
932W2mAakNC3qBybYiKOgFeeliCg8Fz+n/E4pZAfmKspJkLj4hQFA6o0QG84Gt7S9HyyQTY3ODDf
qOHVqDs+fL7zL0C2gHSWz2hn+8QJQNzS+aligxskwAXx3wO0UOT8EMVtz5v8GoNnWbpHwUngJ14Z
u9iSNomJGMpPYpP9E4EeafT493w1PSeK3qcE8w9Rsr/Amhf1/PW2GO60QdowZ2ZhN+qptXeDLBGE
35vw0zuoSW5eqq+T54a30LcZT3vj/boP9at8RAANfb2Q/Ziog88VrT+5WoSEeHiSY8GVXgqGvp93
Epk37YX0UrRjsJDRIxN7O0RboEz2W76+vLCotv6O2wJBtsuWcTrlS4eWQtVLHL78+DPnp0YFYqbl
+0uoUk7TL5QY5diCa+aOZPfeMPAjGwoikt62JbNObF7tmSEXk9sQBC/ON681gegdgAY7XEoWK1k4
63TsGB38FrqeuMYO2n3BAuTz30VebwUcOUTmTxH7Pqb90R/dvEqyxLByCMvJ5a26fM4AjCsKldvN
SYLSu4Xx6VHlwGQEIPNyYPJzo7sPaA36NlQErUAfICYDXfnWdf0KAOdrN/XhUwsCiqmnsjS8qENv
hRcwV8MpEOkoClQzOCK801JYbUI3c8QZrYJGUfG4D6++yyVi8BqngmSVHnwa04Sa9YmJXyJISarL
TG8+QXOmAlh2vM9PaE4riOEob6sxTYKKWxmHgedhiiqm6SZ3dbpNp2z66kmwthMGwFvM8q2YtGu+
oYEszoF2gXGuraaZQg0Vfobz5FjWArcCVRB05+DunJF2ldzBr7eoWu1YRrlylvMClDxQqlxeIp2S
soTb/4cUnau4+otouRqcsCnWO1nHDW7P1/CEHLmwqvrK4CPVEUPf9TwwQBcmQ3N13S99hUUEgz35
11uSkmaHKw+ptT6+F0IlvqCH969YysUS63EpHTAPl2AljFIv0dg26zw88CaS5EfEJ+FQQ3UtOTk9
RKZAqEtPIlQSUFobNA+Akf1vZOka1cFnLuJVX+UQ1RS9Kv4lqvtzGSXPrbgnlPFvzof4VWl36cTt
zo7wD5crAn1RWIB3TLV4X3tmgVfPfRt9Df7XTl9yRtgMbU9ZAOQelXd8msNk/TunByNpHnKVhN/j
JTQOkLBOapJ9Wq4EJkqMu25KDqj/WF5SQSET+c5DN8UM8qy6YYbqiNBFD7s4hGGGlPV35rD5O1Ms
URh5VWdcCu/b77KJUSn1sVK+woL9BZ0F2gYPD7sI5EKrzSmC6uyosQEChKOEQSolNfpzeX+U/TCH
tF4/FHNEC0JQmUFdA751c7IMMLVlr6UiQFfi0r9fyK+M0r5BNUt0LOKP+46yoF37I11y3GzZHukM
axT1dxdYHL2k0/M12MFXx2y2/1SFnmFbjVseakV753/QORc550PjRMbBqMl8ygyViSPLNjIgmuC2
oeeFZu4GqvY8AFitr/t4zfLPoin5WUXXQB7BtoFSZcXD9ypulYRQ1jPAINCX/F4dIog0gQgE26AN
VWX635TIqJXukekrEd8pd0LbEexrm0F0uFo1YWSMP7lSmIbO/QNsFf7lEq7ChBc0und3wfDfuE0D
YsOFTQz91q/MnKoHBwmBbKKeUWZ8/KvgRU1ETjPhHr3p7H+7F4aVja6aubjgng9AcIydgekx6jW/
uiZ6IFplFEF+XD2wJIrvZywhctB0mc1gh7ie7warhGWmZAbCq4AcseqHBoQtb5qQmnMIkvfxTeI6
WuRK3AraErtaVGpdPlI/5sk+e6fR4lSaFF90tZVd7W37ciTCKerVk/t9LGy5G55K3NNG10EZCy/c
Z5XrQsrDCMVEZtc9mf4FztWao+5F5qTg2vOH16eLOJF3l+iMLiFy+R1IerYvLRrZwedA7qSrk1jq
wFGdYhxB4mBaOOPQb35SOUlBsOVZe4SKQyL5JyNFhJtwrBBavw1eyQics8OlusATXIw+usqakp/W
7ewoyUjK+CYDVm4bgGFBCGomhXqEVfiWeNIwdHQVFAWusdIijRf5MT6PqTtnutpyhvpr60+lSwHX
RHa5LJz8GsN1EVJvffLgUnZRcuvK3lKeLDTG0gmsr0Kyok+xCj0+RVbmPJ5GW0OXcxY0OP0DMJ8i
tkYtGr2fYedcctl6QGpjwsldX2VxryHdUp3QNmOYmaMbsSnaQXR4nsPoI8kAWVPbRpvC/yT0JrNX
ftEMk9EpCj3xLPGhiSzoElKDUW3LiCsO7pvcypQWU5/NuXAAV1gdYNjqEPeRdUa4PzBanWo4I7s2
Y+JZeilRu7NfLeuScEf56+FMPK+o2uTcUEL+yQQ45lvskVbSzSFMQTqMJqXCMQyqS3GSvExjJIWb
alO1c0pTbQ+IgUeNGpc2JPeOLqRw91RkfKuFHJ3zdf3YSYbQLjOH5cJLsdPVp0IlDyT8anhQOkc7
42rYNvEG37qYfyaKjJUZ+yvyByTadGJh7/GYnFnpF3DVx16Bpv34vIGfEGS5RoobxDwvs59VCaW1
OPlPu0rTk3Yb8ND+9x1RDIhONhjK2BFy83tRrymUy6Xr0MgiLNJj4g+gi3Ls2Ln1cj5599+5y149
fQMYflqHlwbFDkKjntW26ROnSjQcwrrhxHGpLH8OyGDI+k/aNcFV6G9joXe13S5ISOd4kPVKddZE
qYspBmjxyiUV/GwCyfEh1CZI48imZlwWqciX5/8KYcVkVvsGhP8f3AQUGKnT9rN/TC0L1CGRZ1Fq
/5U6zI+eMquNDATgdb8u8RaOwzJOZ37LXVta2pDWuEMFBBtvjAt4HC9E1hquAa463fK1i/SuIWXZ
UG8XTzZUl9tQv1vo1f7Omk1uQzhv1ofY4T5DknpnGrwcwzbT6tgDMXZYuu9mIMakN4LAS3erR9u0
X2lOGK1TipTf+z4wR7udklgqwI8W7RpG6fMKi/GGGUtIfYoPW05Ba0wBjJvblxJaESoJyQXWoiCh
rLqeM8iTe6VETTBkHzK2o0yL9hWBsZlMwHm75psFHt+vQjfjHy180pzoH0Mf9HSroa9Ma0NB/RIq
qMHaM8HfQA/zuyTFjQ69b5iP0Kpy7yEIBnLGMvXSxsVJxFleQzqG1hUHnpOsn2P/PtAyHjYGXqO8
J47H9m500K7qcpWG/mKtiuJQ1aRRSPrKNLRXyqQbKMUI8oODJuAXCD865++F+yI1WRHw09CiVeK+
YGq3J3Z2mvVn9TDD8AEd3mw0qDJrh8i3UiWzcu4JF5h5tUzaT4Tfua9p9qt2iW49yQc3mHg1Q1QW
/sVNceTqQpVLrp/AqlUhZ1f3nvFfdGqGvHgZ8ToCRoh1pzRKsT5l97Sf6xGUhEleAVk/65UPWQLS
9n3X1N/bBTcmgT5SKKGAWb/mOVzQ0gwdsGbQQt8wiE+dK0a277LPoMdaO6qDBnSgdNUrdhfYys23
TS7HO6gZMYUoML9hTfTK1zd6oc/5NiBl/b/azHlcHOyfJem6SsBGARz/Xo+QAadi0IFUvKoV/LCI
WY0XV2gyqIJSjm7NoR4tg/fSjY6O8v/hUyv3RjvqDP/6R19Y4D6J6goYal+fBmLy7pKv2dRHizQY
9BCFzxamK4ZWUDG8y0wWsjGNglyqQnXT2lo8Vts9ppPiLm2D5CmnAe7+GgIpUcH1NO+0r3t+KypL
/NWaMUrz1ACX315ALgx5QCDjVoBhVZAxVi08FRydc2KTzNRB7n7HV44DIkIoHkr/JPCTprsGOaC2
/PT9sVu6YjHcylZihFPA5TOMSnPilQDBpVFvfCgOve+kCynDr5U0Kw7a43MMnlbSGQR/flZoXStH
Ffrc92riywy+3YNOAVYV5oIRL7qC/meIS0hJtQ8b0WzHz0gszleN/Yin2v9yabj8XTi/r9DIrpBv
OUgfNfPT4Qa4knIrbAN0XApK4u+8WNCS5zDGK+ruakGanY4IMWi/z8G+AiTbVVQA7y//xqTsyg4m
KPGl9RqP7t7J4JnGqrhKLpHvdRDWXf1pQR8cTsbJVu30m3tTmmUjDdRtYyIr4VCfJdTpavfdDDsF
sCcUKRfmy++f1iAg1npOlFeBtsggHQ9s+ji97mGr0YUnXvRPz0EwOGSBIVVh0i0LZCAzU6B9+Zpl
xBlW4odVH3m6WzazIAFO1gPQTRG0WxSPpaRLznrOWSMbtGBywsXBtNmRnusX9Jf0ooqpvp28w0YU
NIn+q7edUxfC/e/NBE7g+fPyqgFGmArFwQS3tkJxh/eaICLTYEnCEKsA+Wy08JQV9QgpYEZVNvev
C+CT99ZGSbKtJbTNWrL0LDA8B2AVrTPZru12qrlnGzslaRs+jOdgDE76DnzNtyFDvKvf49fsCfSf
yZoux9KZUKxTxM1ZT9l6iJ6n/tsGePMiczmX7pRTVMrZA04Na4tzWBOPuJ1SFk9ggW7xr47P9kxO
tuKGdWvS5Al4WIStwdmmWtg3ef0lD7piItLOePDxLV9vDaPcVIR0DZFxhSz/Yx/1hvOICapkAr28
MAf5MBtPi4y+LO97uSq1rM1HUHPz28Xa/SF25u6yaTVURKniGhejxi66Mq0QFomYH04pgCD3NEvD
S68UvU/uhvRR87QwSslBcQFg78RHYO4PXJam0+snZhALfhtmorAupVVVUsyn4Ebxc+d7B5WE5rP9
mwnMwRgCV+Q4ZJMAoYyaUwIxY+dVWTMHBWbvrgMsqush+oDmOiJsc7H5KVS68l21j5HcgkonpfYp
794OlC+UBh8gPnhZitxHVjFH/PD1eB51xpYT6o+kIrZtQt6BTu4gzSrOpiYCteU9G8qN3bujcC7f
edUuGMofekfwB3xu+9p336cmcSmMgSQgs++JtWkFtmz2EPyUBu+fugkSGxtmDROFVmqjm371fiHr
eSLznL/4bEXmRJL/NSx9XWHSHKESmFc9s7UEKXyW2juQ5zMHpU5NKeEu4K6rOfRYKHmvg1xJn8G0
6rds7COS9yuIzISkqYO5LnxKkgvkOwz57yJIkkhAbVLLnHTgsl8uNFlFMEdFHysoXFiK+9sfl8+t
eyvtR73M5mzZbsARWl4pcDYb4EdubkQtVsE+3AB92jy0NX4a7luoqPKT78YrdS+Vpg2i1GViljM1
6mrvK/Jnkosx2Nf637SYpUYfNprX5z6y7X48c19GSFzxfH+OaQLv0eO55m0uqrO7UypxBOTPPfbg
5Jx0YSApHa7983UwZPs5FgWJKEBBprjA//bdR0rcEITVbj9YIxgMZAyIE0JiBkEqQX75FPnH+fIb
kfwJmxhwZD60w2WL+LDda87IKgDbETwd29byO5lu04P+EfUCD+zZhrIDV4keqmRDfvGcJR7Vkf3U
6dpnLz1i+OusFLLL9GsRzEzR1eVbMapP9w+w+eo7mR60F8q0mJ+KSIBm+1pEE9EBPUFvm7Ar4uL2
u+VAERZ8BdaXeryhbJPZepvIcv3jTcKIYiBfDxgFT9Ne0zIC/eru74gxSvTaa6RVJdOHvJpTYeol
lPBRdIZyCJ9G+TXMFZLIqkSi5AbBNCl9jQxsyZDwZvEnhAvUrQQpqLyvwdFLhQHqwAJnzT59Y5eB
pbDvf6HtU64GzYabZFr0+6MIyhyZmB8bnVJ+Z/UgdPNOHchm3ZKalBtF8yeHnruSYQz3DMHEtfcE
rUYF13QWW1BctCXbtJfE2KPnGrXJdmD3RO6NxNu+UQ8ZXqc3v5ytlTPdwsNlMEcE4ibzGTHX2JwM
bYGj6WYDgP/pgvfgcZwBlFqSb3qe9Kp/3Fx3ld0m2/+rSad3GflNnmJwk99x27CNQszXtNyTV+qF
vcobnJSZX+BkHh6xt9Hx3yAfAWSFMFQRxgzGttgFTM2vSQ53oaS5J9a5ASkqdCRThnlXC3WkuGPE
5Dfr53F0Z8HSdUTDuklFmEolrgh7+3M8gdSpGT70rgOx/4ev0tSpK2IkeCJZ2ot624FNu81XK+Z1
gW9SsWpcekwSHx3cg8UWFtenVVBdVsJi85yo4tz7Y97vnweeCSMdJi4RX9FviSORaBwObVWKFiyb
Tqxb7J6L/nbRJmxb8Q0Xmbq+45Fmt6F2pHbXqVgST/yUbPSFpwLeYyUkSQwxdb2fJhV5RV/BxzQG
BGS/02pQKcrh32UsjmFFvOY9pFW7So7r4GgB+HF4XGI3d4DRHWDPketmlV88zFb/tGxcjpynlXVl
w2c0PH+Ng0zXIj/aVwJ8A650lYUgpiAKe/cAQuSF0XHA/z7EbgBL/6sOHsw1WjmYROX9ufkIRhEm
QSMHv1I+VLlIiH/B8yp8qYzbSjQFLdcw4jLnCucG53SFosIa1EVTulLNMZ4aIqbnGTUdvsW60pU0
zrdj336s60biYl4MklkP6lGgk2MZ/X5lg+iSt13UeRgrhRT+OY0a84RztvfhebYuCjONOsc78apU
76o+adqCjWNHfL25uR51WAijh/mqc4v7LJfkpdg8U8wpHydr7uX4946MGecvYJC+HVMh9K6NXW36
YHvT0i2uogzpdF9UbsuV4EZAVy7Cd3dkUUEXe3bExkJ83HrMExss25nuU3mSmmxa8XrGBroB7OUt
kpc3AueMCfs/mcKVmgPwEhSbo9hlibegdeLuMpNP6uESN5ez0sl9GAsKvVL5FS041UaxWaZxOYFm
dJ71BFPYGoJWEgF5nHEV3urh7F2VL9VEjdc1/kpV69U3oZcVwatA7z16wb5hQKhI0u+IhnBeSDkL
vIr5wqupNrtMIiGEoZcPX1wEauXKMWLRtbyk0Qh7YDHmmhjoXyo21uC9ySbfTd4LKlnK155rtBoc
EHwqWPuXlLcx1z/IZgSnS0s6aFgPn6oPN8+tNnKwvVeVIaXJXJ9IHKSEU+kDKQw1Sh/aVywhMVKP
rbLaMkv2R/3/9bhwJKtk+gL3lQDqX2X65WNjW5fPXABe5vPk1ocAIjT0bkDHEbVH1s4ttXAFYJdD
ld+3AmyWnZQnI+fQtmcxXNmQwp/HmcOZo5FkW+mY9NSGtltjML9Ffuq3iZUjxZNlbHpWeKdkfsJs
6aDsjunjac7JKfEgfOJ158dCkTEpleHCYeXrGRs5ctSMRygP9+kE7TC3CWnio2F9UijinG6A3ii+
w4KaSm8KblbuqDgsNgx7qIESYzoNtl9ZCCmh96enaSEbkYd3oveU4bLvEbNlKlp5+hJK9+D8OJo1
veGsvKJiQz99xx7wPoKGJdVkX2YuD+jfzqzn2PueW2qkbNi7d7xiKsX/fdiPSp1fRBWshPcQKrr/
EMbZlitBKxiftPOCSEa3lXZc4Ystt4aUFTpTto4FEZFo2yaz3I5i2dug5/e52GLD681m02HzfreR
7ixUe5ANCn3i33uTsi/AklFPIy2Qx3FICtcNXkNYr6YS8qwSa65xmJZ2mZw7Jq9MRtTZbRW2tsXr
z+YMWn2m+pKTm7pilYX90pkwSHBNmyQIw+5WLL/drALnixzcGUst7yIpoHXbPNypErvL9DULd1u7
dfPcsxLGmYkz3OtOOi+Oy+jFeXcJfyzs136UtHXoxKNbSWfMl4tNuJoRSC4RSliPz2vEkslcB80H
L8+fzMR9HAjbPTV33XYPBJdCru5iiobnjVzOt3aX81faWJ+i2tKPArxhGQg23Hf01Yom/s4puXm7
fpGOXQxvxVb2oPWKUQJE7/P/XUg6P/jbqMHXpRQVo+nr3f1k9DzQNWJDSOI+6t1nkjEfxxsM1Dm9
sceNYYdDU3ZjYjslfeh5DYmWZkEtbUzBFH6iTgJsnZsO82+A1OzbfKvDdTLmzbEt9ME+PkZZAskg
V687ZxFqdInpMNihN+wqPy2itLAhjAkpbNYt5/8UG2B/P7Ut/JAiC8XDOcrFH7b80/U3La7EyzKN
vkvH6YWUTW08zYOiLTL0HVRFyYKVsyUw7HT8eqNvngGJt6NVMOGVwhEMdKcMUZ90Wio77tWm6ERV
9+wYQusZ/xts6W9D+L32uuno0EoKGWG3d6Pldk2Vo/PaieUFPDn3AV5DFApoAfito/xOQKZCK0aR
hjdm1Fuv6QWyw6Udca905TaLgAzMKQLz+sENCiZbf7Jim+7yTu+XLFm/KqBsj/1anH0Zb8DgTsXT
PprlTxDYmeNx65I4CX0aJR3K2BsTyeiWFWWUd2JyHLjVuaYQUdUp9/rL1OlRgqkYRdNyqL1QuR6o
GyfPF8Lop1VLBeEpIvPWZxg+INEbBUMxPf2UvMAMTqEB8T2a9Q9l2rF03szlTrBSffdTHVob8pu3
LOcozQrXUdn51Xn9WZ/493BIdVLDEjyg1hmEj3Devh19n4DxbC2OLT3hZzK6Z97l7m86xPtD6J+w
R4u7LZBzD+HKKHQiYTYCdmvDdlDn5mZlqbknAASD9D9tWfvkHefafGP7wj1OwjI9YAp400Sxyi1u
bHHCHIg7SFDIODDufCuHtBS++2g1jn8apeywBbZJufortvDvEBuw6/RwpRNOc59bc7YU4Ynx2cFx
ZDlvn6iDqrhXsmWzDjXmJpvieOlCOwfMA2xRMUMpgwR1UCpFQCj2ftPW5ZpQyb6gkggpln+ElCpW
EtodNGxrdSDNXB+aBghcgi7KOz2va2PB9kD3ObnnUO2coRQqq5IsOBotADrJo5P7fGhoMS1fXNkL
fXZZO4xq69ziMvC5EDjewVLLKdYcICmqY1Bu8qM+qQ6ETPzraX9u/9Ldh1aTgFaDxeN4xJokN8vy
ENFDt2S3MpTBaEg/oBU1kJBPzNW2KSDZx0oqjWel2xQwh4IDADTaRLgv8n1pBtSsQ0fz0M2TFOk+
kc1wsKO4+uZpUJXwRJIHWTScbs9J8YEcyy7FZvPCJ2BISLcLCyLce/fgIHRUc6apCvD2kr4M+Di4
vFLl5THaRwtcD6pJiiL8nZ0Pab1IEIU4CdMw/6aRef38xmiKzlXZ4rru1D89/zWiQ2JM7kYYmLFm
nGZ2HxOmJWvuC8dmj6WZzjsoDfq9LM6Ah/o5PmPhsYF1UEbtnDTUN45qCV9wvBsc8KihFwO6Y7X9
p+CVSOw+IbodRUb7LH4eoKQ7MexBOOVGAIRj9wGsuHka5X1cS+uSfB84nLJXdSEakjCJy0NeQVqq
2MWE+RGJkvRY0qctq/5EiQlwh2sxjerACc9QXxeF/5LJkG+CzeziLhRhlc+Mty/9btfEUR3r8l5W
aK5QaFaeUcwSOEdqXAMGAGghjZ7ct9y30wWSsnH7/PwSe0gJ2DPouFZob1biw5vmzGcCIXItVx5e
5/eD3lm9qz3O3X6U9TRC/vtaRCE3zjnAWIFSp5oPlo23p9HMzyVdYGr9C1jRjfCCOjFLqXeWQ7ah
jWdRugfU3+vu4osyRVsQCJITNmTSm906DDyDNd6q0Dp+C6Ju6LsC07uX0m6Q++1ZG/ghue+Vlwn8
funOUKfLvYo195hTDBNbmyOO/L6sYUkhV5KHqDpJTrDCN8Bo7AkqFnIds/rDp+rn3q2dQB4M9l4Z
2n468hLL/WIN+8DGSfyjnkpDaI87o2EVkgCGrw7I+zHNTgPW1DAk0THVQjzKW8WcFncXf3xUHmg5
Wot/CKGS883c8wRcFkdME3qIoFDeYlD257yYrnpMOJ/Ei1WgGSHksvxfXzOE7VVcoFpmDHcS2+45
9ZtHGlerCims6W/fMn8NDs0BZBbeg7IMJ2Mkj2oC/nhjcnL+qNvrys8QyTKxONKQ4oJNNkTMvF/W
iWREpSrMQ+j7hf1mncdbFhCHrEXwoDeujYflIT/JW1ncBRbkSgUZbFSpniZlvwxPUELhmiuJryky
9zal7F7JPQGM2YfriebaB/OxbCYwROXlBye1uPKCv6J0bdnGd4367sJH29gcTp+sc2IPmbzK1nIG
vwmtphP7ews7NRG1VY4k4G7gcsqxccDtBbkGhmU7JGClyGX3/LOL/3eH6rqjFuaRnsb3kqPeTgMM
M53FsED1I5K47ID9NNM1a7/QPaqzdrUQysDLjbpPF7EAaduXDCsmz/KnRlQg9WECtcPKxg6tlShh
GTz/aw1Ba8bW4wvDvhwFhOdnS/WbXH3Umge3j8TNX4P8jySoX9eGLtUIQLUvHdKWdOU7Cy1ixIBv
bboHgpGb7rtYW0JEcZWToPmuDeD91UGQT4GyMmj424xdbjbu5W1N2vzxv171D0/jB62OKwXrzTKy
Hl2hrkn5ucpAYkgWvpGBzIfqF36hMUito9Sq1qZ66lqliA5xzZ4rw8Wcnp73Rg7ehBepF8HpwhaQ
mRGwBv8XbwKepx/1oUNfmc43tsdux0DW9CGoWhXuY2rUmESWNSrLPyieEXrbvmZXHjyq87/P5W2k
59LY6TOJcRf2bmrfON+kRcG9cG7SmbfhbTMPOb9BOjjwjiSJUbO+fQyoggq+xjbfyDuUSnnhL1I5
kvUTVb1DKACKCcMDXwp6sw5Z2DqBx2uo1fG8D1+glZFzowyyMaDVaNwrRLr7DBqpgA3op7fcTEr1
AXgDDejjQxaZnbIthAzhwsF1SlsJQQL36QlbuFihD/3biE4Qghyv9cgkSAvGfes8fhksXLHXv+ku
O3GMxP2nYYMKmXPaqQGZsENDeh48ilk1eiXGXO47dfpeKMi1DAa6B/g7ofaNQ0Z4pzB2IyGUja0D
FqTdZYTN9mNt2OmIc5f9nd2DzhlmIoiFyV9a8bYx1nktTBA7hmd4NsaHCZVROdxTovmgr8XOTwus
zt//0HsovpABJ61CDD5RmHt0TA8ljADnN/wSREb4lEI4je+b4SyaRoVfADSdgYBD4o4wCiA+lsp7
/hd0lpepr4hUGkQhm9GyVhk5RUrnAm9+K2Dteqxt0hfY3/36+7QkpfG/7lRZmpwS3n3n7XjMD2Zj
/+IftkHJvolzMA96W3Rx7qd8Kk0+EoPYKBJdgYkUDtdYkqB+wNQGgFTPvhyw5ndseWcbYFXrGSDe
/0h81rPwCK3H66zli4TwoFqoeeUz150CNMecZHGadrX/o5/EOposrZr4XotiFqhfXpeTrkaws5Tx
nnbPjs2mNtoYsv1I05rGwjIRTW82Tj4FkGDUkT4ybgzeHt/q6oGOCAA0O6sPZ7OB44mNju3F/x/H
Es0rRyoyUVuOYOXusDB928ooZ0LFpg1qXxg5SqPoEWHXUg9GfBs3PvxsxasHKSpPjInxMD4hQ1hb
lwV/tdwKlgy5rFiRYZWcHmVAAuoaLpENRPxjoD5jw2+hw+jWxA/ZamHpX1Z0FcEuUN7kIGHZPxL9
fHys6/Go4d4uvNWl+DXHQdlsE8aomR2M85M/A5AA8+6cdPh+gZs3yUK+IlZ016KA0gSadUxZkBI/
fL/ix5GgTjBtoieQGpvzMmGZ0PWHZt/ot8Sbv8P8Ty33lRjc/zajoLznSLH7ftk6Hd9FxEFeH2fR
m7PRD8dkpiajUyYE4Qo+uIflb4DEg4yGWT5J0/U5TTZ3Ctj/X7VnQffAOPwWLvIhQVeB9ytYuUxn
D863qq7vH+5Hmpn1WrtV03h+9UfaBOs8UneN8r28Rfgj+L/Wnl/YAr7RkqFsaAaFZ0Y4+8EGnC5r
I1AM9WE3KSyC5ZrD5GcifVyQZDfyusGmVadtDs74P4ofe4cuFa00vuQLrPDgemuHRjECRA6YvvTE
g+ZWQXMTa4uuFVRd2j66dNj7iSKvccRU8/L2YJ0/Qu+HUKZCBHiTI8mw3i7dxEG2s/bJaBH+57rM
gTa2S3VoiVEqYb0vvXHMNwZxYl5y5o9t7UvQQ/Ntli+5gtHKVKTItyEmfQv0vF3dAqG9Aisz0xsS
EkQmGLBGuLQL4jHe1KGeYk2Nilc1YLLS7PuTurkde8row/SRYyuAMI+rrRltjLW/C4SZxPb/BDhd
eQYzmrrzKlsi2W+QlfuMFtfQgd1EeSln6MLN1u5VmCteCAIA3c3upcba/95Xn52X18HUT6UQvCXs
IEn4X0Nnm7e73/CpAX1K5Qk34jdNRDgct7GUXvMChfrnV2MDqqp/KVY/lMgUZzP1VP+TA9qZYPIw
ohwNVR2HgFT9I0Bgn3VFa2UgLcAcPujQeZgRNoYSwLk2x/9QcZ7n0X5fSWrTdSff9IUoS1xiSffc
5ov7agH7+XFY2Bvkbgb5f5XxlaZtdnmAQggp+PhL+nYtgowF+ebTAIZ9QhCO+JEixsgnkR6lJo0t
JEl8fQYFu7YdX6KF1/JnIlBF6KvJxE6mDG84biK25HT2Hb4s3I16DlA/+3sAnt9RQ0tP4iST2S5y
aX+y/oR7/SWv02FlvRT8UKyNZxOJphAHxHGeCg+8HtSnvEngH8xdSIFulCnopzlhpDMwFbvf8YpX
Jciyh828xjoB9j5y/1QDnxelsmhUOSj3t3XoIoWc4DjMN6zJJaWmuPd9na+xnOsZfZJQas6Z1S9B
fjX1q0X1IxEBgvLeB0EbZNI/ZZRhKofN0iJgn5QO23CmcaXpODtPdUG5estHC3Uni58Eso8Wq6GU
KKCAChzTXAN9I1M82Hajgz90Wt0YAz+u5Y+nROVxLIDTHjM3EU2ZB6x7Xbo/377T4qRLNoQozvyF
7HwbaKjhYSUZbGjReRLyFYf6Gk2yRpwbBiDJ1Gu6Z4CPByfxUtUrQ1QYFmTLQoZNjGLYjONzodj6
7h1uRFydHzsftaAqL5VZG7pWEJL+joDcw/CsgjRUk/tdMXSJLyhZOJb6TH3hGhWAUus41VOA3D8u
1spoTHCPOiNe5+8co7LL0oqyI3LSmHYjJi/4FGtJvXoz8PkEaH0P+hq26zwD0woV6/nPiyuvquI9
rUwS70owYnbqUJreUFC1a+9qFYbYyNTG6BdEL/KzI2b7adWj1YVVgUxeRIrXcgQK6vWBmZQXKQkh
gDaUZgRcnzYakfnC9WYWEJIA9u3x3Fd116OQcjEY+zW9yyhF9B47ky0k0z2g056uW8FqIaaKowyg
5wAX7/8EraHJb86U7mcEmPUT8kFBJLn8dSI+9n8eZclfYAZh9uplUD/mt65oWQBkQiyCDgCpvWnP
FHpaQ2x2lCRY/2dxFWS0av4UJCz8F7OfQr92n4EcxwGycvoMFLujDLKDk9YFmp/kSg7HZhRIqIMD
bKhcoOq8DltrfvrQeT3PoVmoVEM+7dEp2YyGazlXnANfOyrTk7SAP60trnqOQWZdBEiPfCeX6Mow
IzUYxEjo48vV1AXrP30Y9PP6Kp9ZVNyzO0x+dDP3OV12sYy7TpCfp5AhhwDWHzeP6fe9PEmmRaUO
UdYRhyBXiSsW1TxVlotoFL7w3EyArtkaPsJl93SxRn+vUsSERvmCxMyMfqU/ADEBkD1PSrrnj0DZ
iUDbBK0d88VJMWH/6Ia6HKZV+FnGtK+s3WPz+MNU4kI6h0GGQUzY6pg3aUQ9FIooamB8lz+fWBYz
yVzAp4hZ0pKNIYNrj76khOEs6gZfn9KAnzFGokQ7woXVizkLpk1jYFiYnSuQ4m1OOhO3kY/EFQSv
B3F/cKw4oump9NzckFmjtD37fAxmMWcHnfULvQcr83gHEm5AklGKTxrV9kxgEkEHyhGmGDRY7wOh
shOdA8cj+P/YlYfuGO4sgnR+K1gxHR6PKqcxOvy5bwsj5slKDackJwZQNRb0lTDhBd7B61eweXS/
mVwlxmWy+0tqUr/V8CqxZY861N0ksdi7Q19EkkLMOojbELKf4wxNaEcSKmXxh0RV/AOwdHp50isP
XQCB1jNLta95Ot35cIaus3t9DZb4nM4yByYgVjnV+lMqsmJ5DUSGyq5AHJf/QklQUWr6l29qSmOB
hpUqXgHnVwmFozWBPKfD7uzO6kOwVw67ELeC4Vld1NLi/h3kpoehs8etCtMet7ca8cSHlfsN8maw
f6fqSkpWIgxqvsM/C0kFE2U5Mdre3j9wCaK+kZBqUNQwLLwG8w7Qjlj72FYyox4dMgmNDxsUf/b1
XHyq36jsGZ7VtJNIWTYwQoQ8/7iNg/VVvcJNBucf7AmrK1Hf/GD+07YdycroT84UReIFV+KfI5cW
EopgmRX/vH6+0oNyblmKJBqmTBvIeNml0JjREwfRpnbh1yAVWqw84zm5v0ZjLrFHCuhx0tn3+fa4
q/74EzTgW9pKPqmBxY05tic04WneZrbu3SSToU9y3Jj1ehcheDHJsF9PxiTV/JirX5O/OAp+vvlR
GxwKfOJF/ePptqHyX2EKdw1BWUNy4xCNOaQHT9ljMb8BBhYO32gVOSlCJDc6S5Fv1Tqt+lkAx7FJ
qCC1ZXxuNg4FD6Jrhi2vy95OUy55oLZTqxGvImxLmhPWT1aqBL1JBXyxQ+v9FkD4LbZs0f9Yqc24
xgOjhjVfJv0IT9c7uA5qlNED86i5EocNUOHwqXe8yhoFjqH8aZ1pTNisaBlcdAfHNXtuqzDdVtiQ
wAohoL+/lfmk5wZtlFHJYpm6940q33Uw9lEq8Xk1kteH2LjuwxCkCb+AEs3SdMLz/KhGeaR84Lkq
UzzlhpS6tiqMd+UCgZozDNnKu0qy6CelWPcaMmMZKMWsjUGOgi9Oz1pSfD0vYtjeTc59dsFoB1tU
Ubl1R0ApywN/hmkKdWoDAmc9l9HTWXfyrI8HM+Evh9GQUgF+7cKMnvqa7BTsqQmmpzvKebbA+csI
PA+Y6LqkZRlJ4pvPsq0tei51uPgdihWAE0FV1lVzzupJezleLcU7hKEDJEn2OzdLrsG51JHtlL6o
rMP7777sC2Px7cOqiM36aAolGW6Y+P5cINA5ZCJgmA8XKfb1XvgXGLq33souWcESoEgd6oIFMAkK
eT7XIUo4THjOMLLYKRzPw4q6XXkQ8EODB7y/FAztyazNGa0isfv6JxR3qvNyKfR3mOkGMaa72qeU
dZAqQmtr4gwWRZi6/G+WXow5ZvmGqesrW28iiRxo18onU9qcDcOIGMKmBH7xiXkA1awUFy/I6wZh
PlAeq8t+P6zWvswFxUhZqGJzKYp/7qDTUHML/crwjyoEgJHH1G7PEZvMAqDR1hFjLWP5M2xbcIUr
n9K2uyysShY5OZETYfsJ/74lrD1eifBnRuxPh3tuHY3s/Yniry2Xwi7lSy2nOP7zrIe6lb27/YSY
vXGdtjxP1ZBprz1qzlmaBEVnY1a67HTKxERX5zdrQjoRpI1WSmBTN0Q+w+MEEQP4Eyc9kaQNTUUv
ROC1qu6cluglUCKMD+T3Nr2AJre6JG9R354HC921X+7mTVcfY9r/zUTevdJtWu4U/hpldIJeToiQ
FhJAtFjICh9rbybkARP+L+184RuLuO0CahlJe6+Oi49d6JTOaetFzAqcLt6eBuUL30mJFQVdLRm/
IRFv6sXFaPKd6H9aWwt1fyYhrqyBBAzYjoPpAEEQ0nZ2JUkliXJZlt5kJkY0l6G3m5gUlgD/P4nc
OKglAEQENo3xo2zKRO4dx3Q11kJ/6knXfhVxzjbJqAFvbCCrXPw3oDsznug8CQS2SjpwmWobEUdZ
LO5SHg4lH/AnC7QQl8JTY0dplKntQukI6qC/kcaw55OgxqzUpVaedM1L7tG0sAcAZOBL7BlXMnLs
zitDIppPGG01ckzAuKRVDR5q6ze2j9owvSw5YrqTCQxJE0xzXK5w8fVocQ4virXWiE/GCA6Aa+D+
VeH0FoAAn5LRyWt4VrTV7o3mH/A0YRz7HNn2YYoNcFcmJM4DqPVqqHEMiWZifLtD4k6Hp/5A0nOg
ynEUfzBY+5tztYdWhlDIkEj0ErMy+JWCbwWBMUwoqTbUwP8i5L4inwMpUuw7XprxNtWUjs2FKam5
46ZTf52ZmQhJAYeh1ipxWpvraw7A4PA2uopBwUaRjA1KkTw4Es1TXFnxZI4luGbEaEUSMPmcRb/R
WvbHo9wD22ftm7J9BYkbkihE43Pc2omdsld9CsmePMGzFVvXxZ7pt6uUkJ7xtXZ/066wYKij7qwZ
kbktlRQE+xe0z3JzLVEy9CrZsFesHivWhND+InszyYHTWV1VEO/M/TeK5Lt+jGqaCkSLXDCWtXVu
GDznauPQSEf/QAQ/2XcJ+D63esEO/MeQOm07j0/a66AmauyxKNmqzY7gVvkokzD95e+sHx3mLlPb
igKdF3Koqfhydx7U/MnuuyltxyeZDUS/s6jT4DmgmrETv0oXZo/HfnmuPHifRQ8jOc6neyR4twCH
C1AbNDZqz02mHjiw7sxuKWxbVLPQAj1BqE9HjEVWIT9YPTBEdaFMbMh/EfcxL0H97Jrhc9EeVRM/
GUrlkrW2mGEuwEl7hVcwYuRER49psHeGQ+7FuMWQQwWAc8E1O83Nsz1o25pjbJcAN2X7kfX69rLu
Tlksnhky4wdu5P2R2YNJPUpMISTh0sGnt7bH389PWCq6wHkliBiggqy1pVCQl/X5eT83B1O6Cxzi
8ThgyOOhQ8ZjBvBsEMzZ56YrnVMbTqSTQGMt3yEq7tXSrc04s6jM+uEeMbBPhwOoDtlFZ7BH8nSv
ysr+SI3zVUS3cpBSZPLnBk3bzQZ82ySIgVy06eBkQRxFs33OD4Rmrpd/mzB4N3/goGZCcCeveO+H
KiAT+FTagIWRd+kIeai+BzbakIN7zw3i81e+yRMZ1U9KFafojaQEbFGxbfuBFz3BycKyJk3gf3Hr
TP+yG7cKYVvTSzC739hKekn/k60bib6HyqJx2IbOVcaFipGD2ht9QBsSjtSiasMGrw2MofUlPhKE
WkGv3eHnGhFEO60ELmv6oxVkW9OrlcY6drnHDAI+1LHTwbskV/mMEUnvI93iqzRQEIQTXbch7OJ+
G0jrNh6OQEDBpmh6EsmxhJKQLB02kEWaKSL8pd+dLZDaTax8EA04P/gAvZlCQyJL857ztkjafJln
XoAPMENVmNgcPn4811tLLxW+d8+9o6q+et66N/GKgwtuE+eDvx4PYoWv4pwakJIMT8P08FeOEo0V
6p9mgmDWJ87CzVFFkl9QRBhC+a31xzTSj4i+ZNW49a4XF/7+g3fUXdLr3ecQy7DU5t10o+tkzeSe
wAgKmzP2omjhsmdHSL0uL7xymMIb188pPGEy/AtH3ZF+7EUORgnpamnOx6KWP8RurZ7eupSSy2pY
hKbGxv65vs9C7fKp6Iy+yANc16eq0gisj7vNsT/azx2kUkPyBLL5kPYpojScXolajSAQHcb8FkRK
ITLvnRdmCfQlITWB+nY3T48fokYr861+21A+vJgy2z7gD5wXpF1PtGj5s0C4vzxkSX5DJBwPEVii
ekTOF0wVjLSGlLJF/k8XBal+19L/8MCyai0UQ+wBUi38G6gPmmPQXroufPCORc9f9+KTOM5Sd4ao
v2Vy42WbP6iMNH+KxMGCLwpRxkAeLLJn6mu02lqTl5yHC+DmRyew9kepmvLGtQ03AAePfKwIW+N5
PbjEzyof5d6LGMkpBdohX37IAQofDIZamysT+5HSKAkj5XeTpycQ3ywjfHOGnsmCq5b1Vu/P751G
UX0Qnm4pCSyB7xAErgQG148DSd5R4JJnvNWcA87fde45Y+jEFRUD2SqNv2bmEK/WRMS24zS1oLPz
zCfRBYZpSLjKsEkvzzHSWA6ZnXMPGRpNxi2FOD3+g9dQ3wyib+oFhMCD1J/aCWIHzkKc9CBC6/zt
fpsA6X8KewWNnsBecZhsyGlocn8ClDgt8VQ2bSj3LqVcRiDwqhxHq3ULvFRSiwz9zH+aDGiL0RKw
9OnSoV+tYGtDMjBIPfq1Bau0C7lRJ00r0TcXYl7Bc1VqTR7j89TkUfyxkXeGPxQfGCeKOeWw12lo
AaC9qRDqOa48fbZ0OXiEzB9a/vgNJgEi2t9qwr4iW2CJEJ/O0W0WZI90XOocnj9bvwXxCb6ZzMdY
3IEfb3zugKgCew4Qdq/Brmi66VLlrDuPM5allHrxpa4K2GgaSaJFrlh11eahqBg0nBU/42jhB2HO
RgU7IzaTaNQQC3fTM878gZiIMctvV5q2WUUr6ci5SwVIe/4QxpiJcZgZWH/7U6nrGEOIJAV7y+O+
/F2iqHai7Oikoy35L3+5zDQIPEgDXLci5oAY+Vo80WGKqwVCzcCBNdOuB8a95Z6OETwym9tpQo6d
s4RGvPZib7U1NgVv0SKz5Pw5qK0aQRzHnL595X8BGu4A2dv6KgLDXtt5MRQuJga2JGxMeMFNu+1B
+0XfcxoAvJh59RMVZ0KyFfhjhAGzbpgVKW7+a5VVPhZOu4IcmglsMM62E9kr/GdsMSTo77iPy7lX
kwdKfhtLQr7ZRaDJP6o6hqEKtT73m61bXImMVizlhufkLhJyR7aeZysqnV4e9kBDWWgSl0brG1p3
Gbj9rFbPTEjOT7Wy5uJXG76yaDw2aapJL7GsNVWkvlNp7kXx8Ic/iOvhF2KcV2D0NJMbnEd9Bvhn
+PW5yGmUxtdK20GoiN6fieCAU0PELAzMFUhsaIJhj5Tw9v+HUvdP+f8nr1Vbcj5S73otvfnoErqd
XveUPUzjrM/wr3rmGKmhOE+EZxkP4OEPecKoknKFgjt6Pojgd+A6wqKQm7DfS2Bug4fC5/LcRZtk
Qy4kH21j6UqLpbe9b5+e9RSJPLnAekCCC7s3pqk2AtbLFrMrNr9BAmc0+c/g5ZhIDrEHH3sEtLPc
hCcsKj0ejJ+QtPy0AeAJ+nayxl2cW6NkSBlcKOx2/sIj83NNko/xdF6giVsS1YvkpglmOwEqqkmI
jR2VTd3CspM7gOwB9l93lCPpd+K1AnUT09Rqw3ryhWJXd91ecG2Da1hD6fn8J/OAPt6s9KsPckhD
8HG8tW/XSB3eKJRAFChAohvIkbNDyjZ+Z2dQQvSDn28l6i3KYl1BlcldZW2lSXE9KQEStMHdRH6D
2ecvD+z94FBoSk1j6t72Bavn11Z0XtX8FnPiZXEG5UE0wIcCRir09ea4nUo3YpJecFmE68AR5Dow
FlSnIi/iU6RFHeFUuWJKP60oaUvIOBFgWURN1Ki3pZzEqr5ZY2gwv0PFXuc2eUqIgH0RCS6zgWY7
tivkvUKWI4keO0EN550HENpMMuXi9EqjSRMeyRy4/V7zJODy0t/LUwSSQGGd+/P9vH4BFgIB8pHl
8NYsdJPND8vR09M52U4ofmfoxyQz2WtaRXMiqPZDFLFq2FUS6bJQKRsJezILCyUNoCyDK+wLEZJy
y3ZfFi8bCRHaQjhsKKUx4Yo+3dpqlBGCutemGUDJUuvAmGE40Qqa1f/bO22J5za/aJHgmjmK8d05
09pMZShHWZ/5tUGzTL+gYW2Y0pFVXepYWexZulCehjhNFNklM5hYveCy9mknBXDZAvbZaFEUpRsV
WiyWhkiShM3y/6Xyii/B+dib3LSHYhKKb8XyFrOByEwBgOj+Yc6XJaPlr2SHvsPSFUljktEaAnwY
G91MCmDAVSzIEMHyHqesTvw+M3bJ9lVgTD1nwHRqh96QakbMmYwmyfPrCoWtsQR17YNoZa7dVIFt
SeyBeheWqW17umbo3h6FHu12Pn5M6SewBUTp8j9D6DA11Iy6PIQB7WW2AS38M36EpyeOwIwVk8Bt
+k+tFWjhStINHPH1OXzes/Y59UYmAVGwA7XVCGPkTXWPMYVg0yWjKU5oYGutKwcRBbBciHevS3HH
fNkCVHh4/qpyCh6QPUhB4VwfrBUgLdlfFT3fP1FlUi6Zgyv8b3TaIHLrHlP4wajcHOsG+Un0tmhC
qOWcLjBpRvZAz4zxVkYuDQFsJ0rIF0vJWYUY6B/CZv9t4d+PSKj1kXEWuki2vlcCy5Sd1sOzwkU9
iRLe1eJKW8lFQhCtoOoQUvjHU3HQch3eer0vYg+GVNIErPNhI0xDC/yyJQBa0RyyNa6U62Aecwhz
L1EFvSP3zPS+pFv5j8HV9kkSMAw4Eguxj1t0tQQ00WC+D7GUAEn01Z9t2rD/xmw6CMkuiCPaoWrT
/k0WM6+DDYDLrM5c14MlNFn+2it1ivPvO5MvV4VitF8ikKuWy0NgwU4zb38BYwY7t2oNF0GFiQqt
SanLupF7b1j5j0wHNsl06voiH43A8gdwupHqOPgk1j74EoS6lnR0/KorWEQmO7ToWyG62ufzKijN
H+33pge1ZSpxewaw+ogD1RnlLeqgr1KVRayWwIn5w/SFzjgUVywSQZP7+AFV+vqE5V8LmKromEsq
krR45/eyzgTFplPtro5TFD7urXqbNe1KWAnFUOvhl7RRO+HQYvsLdqPicAUSzi19SJOXJAE1Y9kO
pA4EjCjS1HI/uTCGn0BlrvWVYxYAmZA3HXS08xtik2wee+3+/fMvnIeWwBfZ5m8dIfbuDyVDC+AS
ZXC5Mm5v+t7ZzvtIPGicPB1PZaFywhTBIV19sgLLiWrrDEZVb6xXyIg8tu7VlTldNpr9yB8H2DjV
U/yea9qOXMC3lEyaCVKN0HYaTHEbgtGCB9qeUL+lSu7wulpLj0SVS4LZ5qqOb7ONPlWxPYKSCVPO
SiSBRSbWZix0MN3hC3SyImnW3C6LVRFtTwL+dnn/JPXA4kzaqYxJ+B7E/QyYBpoTwZCLZRI4cEwo
7S623v5p4Vt//z2xcMndFOaPdg1NyqJyaugH4nGjC863dNJdnBsSo5VJe0Yzt6OSUJOX6Hv+tg41
S2jPjZZQJ+/CSMTs95qxCpbU8VuIeOdt86w1L2ri8i7gr7V64E+hR70+zZ8yiVkZ7sDk06DpOHnI
25geD6krVOw3nbSWOAWyfNoG3ebnzhG/QM7nu7iId1xwXv4ysBIWl9ps/Zbv41W9oFf3ZrxLkdpI
uqFYHjadzMqG/PAM4/CcB6q131FbRXP8KJN5L+OCtln7zHNY7GvSW0wzn+1YHtyv4SU1wcvlELPd
lH+LtE0GDMSHHBZRveJUSaWUdKskWbPUd03CMp8IzOOq9pGAHCRPC3x677H8JEQjo3UbtVj3qrCC
6XEfZ46jdYfbz2QZxPM1mjqwC3RWasxG7ZohyLzJ2CE23mygmmIxpjks0oMnrkQMPv82JlkSE+Yu
91B3Vb2+8hixfbhldtQc9kOqsMQzoAvoD+Sy1FYNnbIhcF7fBtrY48QpSqvQdvUlCc4wu111wnjB
ARdDaZiQSz/VQj8+dya4apPpgPmmTiPHzL3Ouh1PJHQDcvF1gRTqLXHlO6luaKXNFV3Wxp4mNsI7
XzIE9XcAx5kRbwcHub0Bd49ShEzz/hDKyTmw+PHUNM8pQ9SG/HWWd7yo/dDeVncHNWNrDofC0j2t
O/g3XalkAz9Itbaf4MAUi+W1/3f/CuUTZVKADqqRSQMK5yS+TrydF+w3j0HEEHSD2wD4iNSh2osu
6CjY0Rc3kmjS3punzpHCxUNLsUJ2nx2npz7/OvaybuiTrgjdelQiEKM/ggDnLiySO1lZqXJp1XSO
oPPboWc0rNEeb4n5CYMHpkEL41x2fKI5vWa81ncxlXsbEGs1pgz+Z41xx9hDqKbNKo+QGawrhYp7
WjIwpTRDs3ZOnMrF3cpuEKsLci7LmXxKUMMBMNneZyQB9W1UoXDMWQJJXck0oLD4MYNBkPhUmFjU
BNJHkYLLfeVkJ+0rtlw+du3Gi0/yrxIJhzGpALXl739z/5j7lsFkm11tgk3G7jQODu7IZ3yaAu5G
MJ2R0NxAXzJATq7HpCoFOdutVnogkVs/FV5BdR2bcoHD3Gun69CbMLF09W1cQCRvMEYwzeujYp9M
UX5vKBPX+zBDMJpUvPQ6l4iUcjmMrEvP2lSFlvY8TljWhFyP1XHODFyPngl0DBUH4tBqfWpdPaf7
Mv+/sIpqTV2Oc5TmRc+2NDkXU+JeJT2gvtYnATTNbtNDxeN3EXnUUPuFVZs6eDMWWeT67ypDq+w2
aarpzgvcbaQqA4ely0/nuFbbDWFTyv76u92GqmkdIJOvj58dpVWLoYp31bZphx//tt4RzC2pYJxS
UQZuzWGKK5eTsx5s3fYcRbNNU17Vp29kMRnEn7sq5qo5XdICGKsTOHKMo0WDtWrjHyiy0utJRPkS
1meCSvgFkWbu1AFBx1ZoWQNNUYtj4OCPk6vyCduFgFuFD6NxCcCyaJQTWPky19he9JsKp5hiXOHx
JvSH5dob1o4W9Ie7up5SBxno4MQrAs1U3xHO+NdKStPPZrCFEZjiK+iHXfi1Xr5qORrtwMvJWq5t
z2bNg5vdhajQEz7sk+aamRxP/iOMbptgHRdpMqAZrLgYUGL9ac0tUXog8MzH/61Sm3xCiQuU8Zi3
V6rFMAlabwWRgYlZ3RJBUO7W7GbSbUFkOxu+S20p8QhCvT21+xJ2CTaOLlNaN6/c9gijU3sFeYuE
eBylEVBleQ4JgIRtjs0UGSZuUJrnVysVQrifd5kOKoIDJJ4x5xVtyhI00D6wsiCa7pusZLvpwGtM
Uaw14ieIA3INN8I7X+aEcHR+Fo5OtbaM8PwQYC+U6sH4OOCCUiTs4LZ1RFbiIhw5K9p7d/Dlyi/z
kJvwG/Aq0nUTzOZq2d9tTmOaBJtC+XsRNYfhGWI3oybHegMn96ofR24MVHDjm1uUBcTaoLBnqa0k
P9yyl6lRG0R7b2L18WiUSzJNJQxVB3ARCXuKr0s/h6xHRiSSdmj6QUasOu7VHOJMarFsZYRbWXrN
PJ6zpYAc9Qods7sAwvLMApswre2UiFpXAkdPrC9we53Zz9qp/Jssiy8DROiD0Rkmi0SHJ9pmBOAO
Pi3cwW7ln1wp1MSiYAM+mhL6nV21JPbGDNklwRvz+oDCMv+ID72+t1mz8n71MYvMykfFiEmktHVJ
AdH/ZJNYIZPlmPm16/h2rNHRAU3AUxtVsJjii0VorTr9E9gMjaHeY9aOEkVSau2t3KUe7DRfTfor
jk0G95cHq0fMK/5HQgniiWoFrVUL0dQoZp12dXHFT6R4qroT2WXWvf07FNcPIaWPP07l501ZqFt7
UM6iTCHRSJylz2Ip2evTv7AkNLOhAL4j5k72nYLChFjlkseLfplvaRwjvPmVw/jdu6iDCag26OLG
/yNSgio/HhEm4dwtNybOHmqXtHYGxJbxQLmHaskpjRVDPSYK0IHfCbK7qFgmYl0XN+0lr06rQwvq
Fj0WzMTWnNlE67n1z5C9nLVqzYZyihi1/SvXPgEKvEOq7FRysXxQH/KYSQ66UavJt2Y2Q7Fj5/xH
Evb68e1WrlR/wgez42QFtmzWbMpLoqYxUaQ/6v8CSr8UHAyFVvmgfurdQmLz9qHAArMDwV0ObXRV
N3+7zeH7EJlyX9XaLb5m4URXwvX5XQ6P+hcVZIABBFQ1B9sXywBc3fN2USQpJdj9XgLuLJILgEJ0
5uZr8VNou8I/QKou7jXfbO82EUCJhmrNtW3eq0Zr4htOk7JbvPNHpojjyNNIZWu9+m9Gx357+So0
erJuhxDTrDcIKmPXuwaKympa0yZsgV/31+D/6oWbLkUW0W0FxrIPWu/7k5TYyTMeJq3TSXd398vy
TV6vS6vLM/gJuIsoaNzUfpjoYHgcV/ane5FX2TV8Az14o1rHULuSeYkajMVoNppKSiU5xZDVs4TI
+Flx0/X/kT0RtVu0cWd0LCxoQsHkwgYz9jnI3XH+6Uzxv4drGkhEiW/Lbt8cnPfuQA9J0VJVSuCB
v7tiUdSKxNO/lL36bIOQ62LJqpX93unBuOd29GsFK1lS51ugGO30a0SW7qS8Z8DEtm1IT9lDWgcU
2XhgAqL17aufDCggLSGHxenx5kFRAx+J9TWg7O2CVqMfMzrpnj/nymku2je0+qP+kUXdM6ejt3Rf
Sgj+KMr7fETj+NzbVzde8pv3hv/SnnkSAzOZpPNQMQR9+gOAdu7aT19T6Z84YA6acRGpxz30/Ec0
E0tuhqafHlglNXxU9zrim6BWZVeLYJPctcFh+UfSlbt/2OPxPj19Fauo/gwTOaa6VJ73QCi8lPx8
mGJmiY4hTthoxcz3wW8A03gCyuolJ5eAgYVBYJkUrZleH7URnwwtQQthGSxb90x4ob14h1BAqzqF
nuOV/JGWhlaYm0aExH0ystmLu00JjnQJStiw0GDWmBzXGag7RG8kUQujr4nfEs5qpCMEo70J7rPb
Blub/m92VfIjGsk6sMuXVSNKJfNK/MbJAAudEsiCEePb2fuDCoiPaparo4E1d7MA37I2/jbqPpPf
aXJlijbrOQBTeUJpS0dATu425AQEDAbFk90oIt12OzZSFBDAdblfBTRW9jkffhMo/RlFE9fJ5jc9
Fgi8AeV/l3tABnT+gN2z/E8I7MTzE3WYCmcFIahScERAZxwjpuIFx/9e1LafO63QAt9J6NPaM+TS
KpYO1mCid3u5OtNThCVcKAfUEyjsFZK3Jd8ytmwCZ/3fsm7FKQBV29m5MElMCvNPpEcKmg3sdYMG
+QcIN/Z/wFQLU2gmG3WJe0FLHWkZk81VuxCpMubH2T4pnYYkM26R0bbVIWKB3MONou8iBQ3earz+
TnEguO7rGTdFWfgBlNdVrCFMxyuH1zzL2Iq7ObE3CLo4dq39aiwVKkWagbgAtFnt7YlGcOVLSxp8
+mg5W/iv76xnu/g4j15w9lpv4v/qmy6OHu6lxZQmdcDod+4Ux95tHpFBwL0nAnKI9Lz8BNYLXY1T
tkqRiNGZlZMbFZcBTedYaj/tyMZGmz8/sd/7skHfM5sL3QOosHPrH9AevEybjdLwjb0/C6eiFqG2
8cDoP8vMZeg4e9D/31XQ10r1v2YRKfxdfJOwX+ZcuEqgg4Oknn9/qtfyv4bQUomE4RGwo//wAuO7
5ia7cESw8hOm4dtN3pwqyLZ7EXaOs1D8qUJ9ujILrj2S8OJqnEPTaA1LMuhrEtnJDyxpjwfU2SBK
TkEGX4cSamRvyT3ANdAFectONqOFHfFdN854Z0jbi+FYnTgoJJfsxWlUyGyADFp8PCAlV2mVRM9I
sC1+ProDtWirluUtqxMKnuS0jTyyNLvzWmILKOKHlDLIcX0oCWzTNNdIAPtw92Nb8AFJ4tyHNsfG
Pfk7Zs4Y1Q0yuA3jGf4t7qyjHYdUjw2rcbAtln6lQCcawwl2jtPEatHeireWMmTx/nJRPRHkmth7
vB+pRUPQGCuPh40X/aUTPjXhwldcyxE4gCmr2UYzkpEike4Mt0Q0Wf6WVIPoxOI/hlW+DjZFo7Bk
1zYIT4MwlexYktm3u1em5/qvbBNUv8OBrkn6MB9j8wWX3K21lD4Hylx96xQeFyrcS+r4HzSeIlam
xRUJdI1eO0KK6Oo1GZiuJDDB5FzILWk8MVff8ANSpOlxIDWBvyAGwUrXTzde+eTLDAi3/4Lw7H4+
38cMQd8GN1aD9IY2Ej8eUlAdnUyCfPUraHJF5YfxLhYl3OI7/McCXUVf9xrft49qJMwXwdKYxujH
kq6elSW6IUw4nOEuW37oWOgt+nyG8HK2DXDNSUIPlmlcUFXRw9gy3Eph3Vtv2AQduLXrorMSaD0k
WWkNh/DeiYCsWNkKiflorsMo9elcREZYFPUml1cUhe9rwINVgLZu+sI4/TWPb78afBWH3erfhn8o
iF7EHylHA+odI6LtzwmMxDAHp0i5lCTtL2MjMH4hXC4fLg4paepM2QamzdgMTjBDHTRuvChgiCC3
QH6dOfNUpQUCwfcXOcLs/3Og/uawP7yiLc7fSVrUXC+794vliRWQe/KWK75atc+siFyYsjfUwQDd
PmJpXp40zA1dDxGeJo+XQ1p2AyNh6yBhl9qmjvuxijGxkLe434QJmBv8ll9ewYk7LEq1HrTDfgcC
xlEafzeIaMODbJJ6Csv8W+QYyw6DWU7J7/4V1ePD03KCEWfCFH+6AQnX8OUu9GRq/sBB24ZqgfEY
qQ0cDNL9vnf7e+bHLA0iBRUqHmbJlpMX20sx5JRDf1PD0bSklnLjmmPCWXpK3FPWxiX9xpP/aTfB
cHj94IDVa8iLuqdLC18Re+g4jFqcs9a1Kty/6cIqHHJgkRskVx4TGIWtZyLYymVXqHCKdYNAVVfE
kdfv7Jxj/BSbT794BqaoCCvd4h9LlNBDniNcXgkvvlklLbQNm+YdOkPCxWGIxYXy4sDVmZTKonjB
cm3AlK77L5aocWxHHxxuJ4NzTpuQNUkTkta9ViRKbQ2lGksSerMVp0NvLBUbrcF0qRSJ8ZzHZa3X
kny9vNdrfN3tbhVLhPTpKIRzxYZabKoNn/wu2IM0cosPaoAoYIdEk1ZLi8e71cSpVnQ+oXbSoWSR
c3+bJ5UptfVmA7oFY/D5hpC+zqLs17lcF75OiakEtgXiqcGO9UQA4Lyer5Qo/iR15VFW3K8mXEGm
8HztOYpPImRoEKI37BKcJ3ispRPussTVLIh4f0bUbO08+rWr6hAu9Bb2s1XGuWKk9zVn8BamJ3a+
z2zVfb/bI5SyWMfK9jNHv0jD7aImX/dFFRnFN421UQKRZetPEGQ72OK+5JoYi2M1tDN/Q2nkOE4T
F82yA/cQ/X7tnKb+/Jet0R0J3zn6mVKnLKZf9iN9i3KR6EYLm4iEiN6l+rbG1MbTXkDWEvozaCu+
rH1uYSgGObCr3xwb/1nmitMM8vnkKXk2pNhi0VRmTJ73mjfJ3+kfb1t3UHCZCNSggD+XhFkLBOl5
KnByagXY+EyMrcu7bR+vWHzXTWawZsBv2LXA+ViD7Q9NSORFiNReNbRHbps4jBDOWLnwWPNYveQc
iS7eAnq1Df3D4Y7F+HdPq/kosk5qnRGdDNTOLsGjlT8VTVtvC/uqP06BqZicJU7oaOj925cDIjyx
GWsth60d+ARGrhNKtPtbwSphDBA/ryK9Mw63TMm69FXyVPqb90M9beGs9zlw0jl1ZwEYATLsfGBh
SLOWhgCg9ntOwJN24lUhT+Ovz/I8fXoSZZu/whgvQxulEVE5R8vpDzyuiJS6HkAII8MLaNDRPI7J
JwGCRcvg8yXv7s6U/jfGfUnFmQeBqCxhd5BWhbVr5l4bBumbo3/qP3syOAhY3n6/IEGMhIvblAl6
jxjEq7F8qEx1W6OJsxPOxAv/l1Vjd+MN3D2MV2QWrzEXKMbuNneRE0ARda02Nm4CeVGaTNpUoNI4
TZfeg8w014w9VF6lhp/xloXVBs0zQjSmTPYPh/+usq5qr8l9nsOOndUXiswJrSR16dGivKbeH7JJ
A+7pXceSbxHQIDXXxrcVfMr5SOOJPTMNLctW7qiRtFEve8gOiU6p7EqbcbOGFa8cJ9LB2JD7iTEG
3ODitirmITnu6NSX7ZNgIKffTtiA4ns3oE77Ui5mzc/dKr7xbi1v/pT3/KKZIE5YCIRS3XcY3FR9
Bq6YxJcF8+3oAV/LTimxryzDZZ5rjZqk4lCnrmEcAt7w2OtbW7ctpaxy6A6S90nMxWOn8cGNw/Rq
x9g/8BHF88REAI51gDOvy7aICZLQLvgrnQImPJrX57wnsl06MWkn1ZLqsWo0dSYuIYLopnRhHCDp
zTU1oCcTJPsx5CiczMR2W0H7oDcu7XlYS5WS29Jk23OkZX4z4cgjEw6+wBhPimSOKogNAOHHmMKT
PU9NJXZH1ZHZ121mElc9CqI+mOv4oFWsoAUl7FBWEpsDiBEQixX1O3oVbLVt+/TJnWV3IH1nig90
Ig6c+91FWGrrpsxR070Ab98bRrXZXjzanvqGdfzZ1bEA02Ekiisw+NfFfvzUSZWFDaQg9AuiBOaR
iX6S6xUiSakxjCDiNfueWDBttwkv6S+7vb1ECsp4Mcys6egVgiUwbO4viwI3hHNLuS6CEGQJmzIv
Vp0P51uwPqOzJBhJW3M/1RonaWnWrvw33UIZ3T+9+nyGBBdITCl5w0t+W2BMPbT6XnNDqGK3Twml
sFZknKBqjxCxwQRgkzHE+rZOJgDWG24U7VW6kTwvfaOAFjrGpCfKQNIApD24pH1KpOD1CYI1I6q4
pPEJkHIVYpa6zKxYe1gE/SkZSzkxk9mZIjCBHYZoCCePf5XaeWk9abKoYgFpMaT6k0cV88Cu9uYT
nvqBhMGHEgjk9rle0NmHN3xUa4Qxx5QeZBSWjWlSdTrfI2YGNRpo7XosbbpCZkhqGjKCAUv2rcTl
muEHntVHXGmXpmJKootBzHAkpYuXbt2g69ru8bzr+ZxCnGcRdPPcuxPPv8os3CCiu/oXcMGayo8W
Y238dRgoTxxz5AD3oEV1t5TyLa15w5mG671beCrQajVFY/9C3rA76mFuelvMGJYGgUrNRHjHmJma
uJnj12CdnEYDbizLOgVQ17ufaR1XrsoLUfT5UMXHYQdh5iYAfHnZHtUKL4WkcNohoyAukJA4pJfQ
PdAp3aBv0daQj32N3F583zv2z3hSqj5whSjshsq/s0AF4nihW67JXWd2sggAuGnjGt9vj7Wu0WA4
Ai8Gc9suYphboKhIxcZGQlMVjxWwWoxyWZ4zKzXG/mTVIhN6KqpEWLmRSBBum8Eh+rjx7MgDXdJB
DvbKv7GpCMNOMrqTbmlKd6L2zk44jypZKCcoDZo/qMcdCvA7heLw23s7qAk5i6diATSfal2CFENi
v3sPSCs2rQ2+C9uuiQH8HL0FbqqgJFz2eq5uQVMKSKQjd4uGJin6BZEzNqfAd46PThLFsZGYOqv7
uY49LVm9alFCRSh+PsgbTX8YJ4yR3GLIjLZM4B1DHUyIpljKiKso5H0ma2k6ODn+wm/aDX0yr1OH
NdxzLOgTu598BD9wBRn8Ltglkhzm1iCaXLlPT9b2h+kjPeiQPmHP3tPkRFDSWUHZDt3J5TJ6PRdS
eky7c4F71SvYzGTsjIKPI2CasJJqYQan8EWziNa+wE71iUM+KHX5rbEqlPZEEKyWqCl5vF12VXay
4uta9AlgpVOMo8JMOt+ZtbIvmMEI5kQcijAeVM6YQyvECzLkTFKVT/1uqSl6lh+8K5ns4ZDL1QSi
Wag0RLfw2H8RfVblw/vEM/L+lLOCN+igoEX3x/yuUVIT9yiu18tX7DA6fLmv6LtMXhlDWY7/Ylqm
BZCWsUJsAUslr5tYphEPxP2Tc2i+w5RFpQ4DVvJJxPnSuRvVL5IlKp87r8eOyFXgifBRa9qgBzYT
Rg32FYGYqdGsz/edsVoyrKxf7mBelbKCXapquE21Mlvay4p6r0ubdijznPp5sKilMxq6TWTsQvvI
XuN6ja9y6JfcXVZAaHP1t7AXOjQ0uCSi3UPpHkdYsVgG4j3PYZPdLPQNK7VVMD4LLXw6UQ5WcR1u
wRh8e6dKk+dQ0Jlstw/k/VwznD/tl7wIMZn3+HeXF+iLhgvhqbHPcJzSxgPmzKk5gNtO9Vd+hy4j
60jhZ76Pp18yysSafkRct0u84vfS142S/uNlr7DNLxrqeQML45wQpudDVKFPm/g5IX2ErZxWH0L+
RioFQAx1iG+7ZbTACnvZ0RpWiAp7ZeD3cENO86dkwzlx0/Qngz4ek2iag94/fdh5FePtIT7SaUS2
FyIieIN0z2UnQmnMC4L703R0ZgwgW+yT4dZMEepmG+vukfifJ1WZpkGcqo4MPm2eSjy49YZT6psE
QNyth3SA760KEIi5X328Xw23+moSs5DtCywkNXK08eEiYTHUrnPi+OFSx8mwsLKO56i8CYJ1R79A
exlAs9MItfLLBrIbYR/fAeiPyE9A9iEQBAESki1NjEV02xzy32+CSw1B+Zba1Bw6gHAD+r8/+Kbs
4Nhzbl38UimhV8lI8VubioSQR5P2ITtReZlF/r+fYmFEGO9j6ecf9IMdxk/lE++rjFNk+ntDyX7z
FiWv1eDeEaqi3YDrZLnZ9VR0z01nRbfJ/n4gx/7yb3v8QW+QLPJxhb+0NcnPyW4USRBUZS50+mj9
b6a5p+uUhHrbQZF0BxZAdxokveWLvquaPu3d+G01R3e1+5lNtybf8iGHToHJGFGlajASdtQyPC2E
JNorirmQK0FCPa/m/LfDbb/VU6LN5bXIJ8dFVwdJoeNLQBeO29uW196SSN0gUKHUPwYrYkflO8P4
YT8lUKMxUdy2UjA6gj+Zf8Fmnq/CfRoI5I/b7UjVzKAD4NjYFKKmmUBbNpOd4NlAV0DRRnkmqEMr
v8+dPK54VLPF0zwFai6CAgKwAqq/jWlZVdWxVaFV6Me1bMh60EG2nQn4WaHRoj8x1nNJE/a+I4HJ
e5zyI34Xu1NcfOeG8FoeuLcL4KeDGsM+KV5GCaRFeg24SpG4vH1eVfrIJ39OF//ZMQ7NNM3xacKH
E2KdLRsPtlXime+Od3rqmptbzg/58IYnBBSuMYz+lrzWMBKtbKvj69ZLgBi7bQvwrU/p6UgWFz5A
LcAHg2486hD8o59/9kRjUEPMlKylsKGvHuYAQQOM91dOVQq2fp0Bfyb32duzcLU/hdoYFAeUZPPf
G9A87tagWYFXzCq0/NnhMkCmq8jV+0c5mZw3kdlc1rQ5u6VMSoncmZMvDQ0wRfdvR1MPzzx+zzTA
RllzEGBVqttMQsAaynm4b+1NsW2igxCjDYEg9Vz/NP2PqEl4vE+jzM58PWMjC4EJB0ZUdTHGOpU+
ix67lX+1yo3qOFkd1mw5cE4Txujl2Gkdz7NsOT3DbJHBPbki95sQT9IC7jc7f3FVqrJGkpmexNGr
zbmNSVU/Ho8pFUYtqZqCwIVcUcmv05CbaLE8oJczdJy6nRjOIFDs4O5Dy3upwh35rZKqQ9AJcA11
Y6H15NtmVC63Q1NWqOVxCoiS5z7XG+E8MJgfqgOGSD/stnTjpz9hJ7JlasZs0o4pCbBg9L5dT/6h
9UhLPxsXAFopoYfPjmpvSoD5xm9Ds6kuodoiLOCG3q3FeHtwSJxiaGybMr4hUa+zRTtZGxXqZrYs
k5vKClkRqYpJRrKa+Oq4JGb73+gL9vVOiSTOZmBqh4wEZO6GkVKoiGcJm/seumvQR1XCu9KLlsf0
O7jmv4O6zCpp+106k+PhZ8Vs8M/KwLoFjdLQf/tnLDMszvfNkE1lXbOPfj1P2yqEeqqp9MchhT3T
0Ya+dQEftI8raFrPy1v1kEel8ovFU6mnnnZquyJg11YdAbBG3gNWHef6v3d3JeGSBOiq9F6tiK92
WTu4hbto7h174q9/ptZ61lWcxy0PCbDW+vQurmDVcvTos0cvVOE8L92/WkclA689cFGY/pD4QsiA
NTDspNvnu4CmEjplA3FHbpjhtvX8NA9Gi2aJH7Sp8WeLtbq/kYCLTJeY4XVLRB1K6yKIu8Xd6XAR
zx3YtDgaV1yKrRnse+nDWmhxlkVegkGz/IAAr7xGJMnaeZOjU4aNF5/t0zmvNePiKLLBUp4QFGRP
zRZgUZzrOWjH3xWkHdiz+3HAjY6OZPhduDVEWEjkbKwR6hWLVK+htpzm1+S7FkGxBc3nBHEGZ24Z
UTWtjt7un/nSHdcWo82DOY7jnKhPBwkC4H6XnYa8ilsiVlNRTZMRA6Lnmo5AiPHgQD3bU3jGY13e
JhcUAJ9+F4urgYuF9n6htHN1NTz0HrbQwbkR/ozQ5TcDyBH+9ceVL85E97gpQ/o7jzwCNEvZ4vp1
vtgZ/R+CuPtgcFfBV+KQCAgNtmire4PZ9l8y3Aj3/7Kic2+EWPX5SyxBRY58U74L6EHXnJdN3NqF
LVrgArq9xrd/bqXXZoz4bp9Udzql1fejSeo6U0R/TTNbvftBzDpLJ94x2h/ojCVUYWZxQ5WicjJR
ga6EdBZRgItz0GcQgS++0/Mr6q2moD2l+P2hr1rvV0Hd+toqXPhtffByV6RWt8ZpHnTJtguTorWM
u0mDND0VnMDkxxMc+lu1ofNe5buBbzMJwAcJ9FuQZt/sX5QIIZ+f5YBxXhkPSUaVJhY32PdhDANi
P/Es9YsUTefoA4vgbNc7cPhryK3pF1eFQvJFKen1Uo8DE1b+2lLFTiIxuChSu3dkk1hqiOiMAgL3
UDNR9L4Q68d+pbPRNxgPCoiAssY3P5MV2gYyTjPpAJj711DnARtjIBWCfS8fGtfXZP4TT0Hfpo9s
bRPgM1P4mNklvrs2FTkSd24Mbh7WZZplw4+0A7flVhrZxhF5XLQCPPw0Lmyg051UPiqolGze9Ola
2Pw4sFyd7Q1YHFhAV/AMKCxSy+UabTGgxM/PTW6NU6pRe2sp26A62lJC0rmhhLyNlQa9+w/q6SQ/
84YaE9Obuz/eV5ToBOdrUVlGrMEEMv1eMigy3H5TMqio276W5iWDLNGcvgi71ktjMOd1Fg1ISXUF
4m/mV52VQ20CNUkI8lfCKqae716yAzzuxllVgiy993QXszNTVpy8uG1sWr8vMPP2lrgQ0wMqwZf3
/BaqTwDtNaSNmMJLp00LfDioAml54cVoUQl8loADqFSzzL2cIeCcxoSkjTnd+/o14mpk0NWCTd6p
Quua1pMHMtxNLL/v17o8Jco3LYigrePcCOHH1XdvDQ5+u2HVNF0V5iunqLahk6AeL2qazB8fCFfn
7ePtUh69EbjeN/QH4dwuOHvny4xfHfbir6yDW3si7JXB3NV3/Tt2Fx+gjKYMfZPBzrxyLfDnu9d6
daThAxCX1CcF1DIxIZY+5VOCltVlb1IFc31yiiaFb64iGG6ZdGd01X6S5AaihxymBJkvXMzD5IAL
mmPQ7Px9wEINk0aw19Bt5DBLAZFQjk7iwmEdHKB7rU3pXCDXUp26f5Dluxi/X8ZL3+01FWMOLAFP
su6zZ9GdKu9gofBZogROU/qQ3yJA8TXiGCqpUpd+89zQZ4s6rVrYt/0nJmP+NDy0OZVt7YR36AZK
PoP4FjbFW7NbwNG6q0inwC9ZSfypADOi2RKi1Tgp1bnSno2PFGedOzAmmPnoQp+htoXkr1V/ghs7
hI5lHv7h/ShLptSAVSQUk0SEs++6ML2kbVp66F0tJWbGwhtUqvp/etHhRIcOM9KElT75PWbqxwMs
SS4ksOAqt0VVO23AYqZzSYXsCLWSoR6ZSDmbm1xzNfvzwhVH5KLHX0NVnV2H/8MtBlwUXV2L9e2h
pKa5xYZfbXK2BtbwkuJZWR29yYk28CG3Hxn8yGEmsaLZMrEz3zF5xlB3to0iS5jW8KEgLHsOpn9u
j1DAvKd2UjTkfJlch83zVDZwI6zcf4oYNYWWJuZas1ePAdfdzwx+UB35aWM4JfuNGzRp4sZtha/x
pPHYtE/5FvBciTlLNgWKDcGzZ4wyXp8HKGAC14SJNs24T2QO9ojCxBMrQpxgBm7apvVD0/r4ipOp
yH2r2bscQ670gZXaUbkC7KpAKsIGc9rJjvVcU3ZCHHooI5yynQkDvTyDMN+qjsiRjl+lLPwopgwP
QlCP5Rykv6QpPHW1Sd+9iuhPp5ccoyCIA0NpZU03vn0AdGtxn3yLlbohQHvVJeWTUHWsJOF5g+cb
WlLA5ym/FIQcLxq5rHDNDubddCeVTPN4AGq6PoOwPNU2eCNqyiZ7SbKGDTfF00Jx5nMgcY1CT2LG
b8GPZnIubuwoBa4nIBS6XSlADq1xxGCkuZbmiqNxIOr+ROb8I3QsQxehI5k2ZI2WXiDCH8KhjCuV
rT6xC3BIPYL4WUodFCoRp9Y+GOAfXeL+MfZAPYfEoRFF5jRoL7cQsc9QUnsKZxqBwM8zjLIAikKb
3okkD6kKPau06BHvmqKwbvjOGuYTNqx8mYk+LoxKUPCBL6aSoZk8O1Jd5+zpKyl9cjCEJg0qT94K
DKFSy4HGBg8EBbx11HGCwT+FUDWVTRz+I7JkgD0rS2VbqEhWYbHdJYCsC5uDIEtsP6d549ME9z9P
rFb9LK0GOv35Tnnk/B3hBIc7JtnFger3cYuw8Pf9gEG1UIiirfXSQm37Hb1O50xVWNU2mhq7iDIf
P+DMs+DtDDzhs9zlrcnhLHBJmrUWDjxaVMKphFgx0130bcpBywFQVuZ7QGgTKx77P1wHI2QwWp+y
ljGU2DvxHVr/COaXyqrUTZyHDaaIzWPZZC2hXz47S4iQAhYitFQWvYld2D4HKWRkJZWK4BYmdgPo
J6leoqR0BznYk6I4Yq+xUKutc5sQTGlvrl96Sm20CA/ZLUVPWWt5pgtcgpkDyM2BODGuzdjnqL5p
7STUC+HTgXX3rMSZgOfTKooBO95urVkhXLmdklrRXKyvOZXakMk668xhvNL7aNIQYWKa67rdK+ko
mmCF0XxquqDdVW7ueGMqD23KxWdbuTvpexPLYBLI1bpmzMPEWHIrHHl7omq/wQW/M7HiF19HrCub
b5v/u/F5nz9cSKyq/xHMgPDnp0u7uBTqEiQxMdZoiHOx2y6jc/f5L8p4AgnUu+169ZtMT2Jt57KB
fSjGONvXzG3JS1COh360GhIlOgVBgdtxTjqAjaGnhZIzXbnFVKOknR0a8cvThLZpcHNhyywyZuAV
MvPEoMAFZeyEWnoq/YK8q2zWRbYpqi4jGT/sjdPV5SOjimUlv+DP3SI2W4h9+q5vl47o2BegR9Oe
pg9zSHSDxSyewro6uJh/+VDQ33TpRalQQ2fcSavhpFzgG6EtbGR76uO30l5jLE7UFZxAb1+TrAtw
w+r7tppsyC/FS7JiNDVU8GXNRSacgn+HvPwNFsXGSb4nHGEwCdmqj0cfZdfn1PoNMNI7FfIt4izO
ucpl7hwvA6DmdhFbSgDTA3W3ZdNe3+1427zhY7lJlFDZimyw/J4dYsfoM1hkH2VZUrNODy4SY06/
NojvxTELhi4h/HRKuZz5krQP85DptTM2NkXj21hmIP72yJLjNX+GbBPvLk8AMvbjIhwHHVymWDsj
blnjrSAR9zqsdAwiFZrziO7XWarYBIOVmmv2HyUZvIPjs1BugO4t8qLkSAvBMsRqcxhtVcELBKX2
tXwjjmJH7homzz+60obbeUqeQEfc47mQy+6gR47X5lD6fdPXdF7uNNFiuORdICBpGjE85LpDcXIy
o9gPkUeENKAuX+0vnYIU7aMU7H0mIuDQgInofjgZ4p+asY8HMawYpxjhsSBQfdM9lDAwu1MTb0lj
pATPJhlWZJUoJUcc9hGWawygUeDTHj2odGhp+vQuojZjlenxyL1upxnimCoH/bZRmKMarraiYP+d
FUI/cpaaoHnS2uSbIK9rXQ2jYTDi7a3skga1TcC+5eH20JPC07entZNn5vsB6e5L0csfhfmYzGoY
budZKZT5Ntb6qL3G1xLFGiOdl9nISTU8SBOIfUE++t+aBEBGycIKFFUASnNLOxHUcJfcM+qz/Mht
KCrStF2waoxLdag/QhyGBphmEVTk5CR0WYkdpBxEYfrorvrklzFarn8bUw2Yoc1pAiGJFdSXGiTz
ZKdo7xKIpvNUi8+kL2ke9W/qxXJbEWF4mpH+0BVV+eKg0gIKapxGcUZwIBU3kWRzYT+RKk6519FE
YkE1WISPUG9WQXtraOeZoauneM/2CfR0Dj2jXF5V+Rwbjh5ndt2QBQ+AFK1ZOik1dDyjdjaTY26O
da8+kgrQf8GuKPBV6yg8MyVh4Jg/JkKvtgG8x8jd9ZC+UefJYhvB6SoefbE35O8VXoP0wo/4qlMS
R5mWcJpH1Jg5E97EaUHwV9hgVqgisFQPciqfQ8iBg0CE3EI5T5WRHXPug/oBXxsY37d2m+jCgZQm
AiV7yw92fJ6AL7wtW91p54iTLq33xs6puxUqNfEEtyRWSrIAhtIRjmEQG3suYigzcjSZfkJGO1Ew
YjPK31pm5GTnfdcVlytnR/o+C2oE/z2J5+HttCmeRqzglMg+XDTk2jlu1jFmKzWylIMe0hM+HCCt
BSQePSPi2/F1fyeffeuGihsnKUelS5vvkjmqxkd6UxOq7sL2CP9AEaojdRjtYPtPiI4QeJ4KfPU+
SFlULE5IkoDDHYP1UyG2j6LkZCItHc1HqUu+x2gAxYcih8ZU651RiK/3i9odan9rJfiRnW/1omE+
dY1k746e0UlQv8JBmm7JCkwugXq1006r3SmlZeuaUJYFNvUah3PrMUinFTtWswQu6G6eOwdXlqgJ
mSvu5oqv6dy8i+4n1lL9iKPG+1b/0ayssVhzst+i3V172sgyZzZvb9u1OiQmVLhIWGwX7vaoGLdg
pK//aL6IyDNXdYrSCkP1vbAyKv8sbo+9AeQ8NjwHQlaR7PA1VbCA8B17TuL4PNZRBDqGdZxEYtAd
q3kN1B1U0OPop2Z0RxYcQd2372x/MxA6uNIx3vDjY91SMyT6KNq8OaUNOwsQN9jaM67+zbDE8yu/
zlU7dU9SPkLR2OnIAmWjoqkf34bZK0otFtWX/l7VRkRVAtqUVoGFYghtzsyMlSkmsun6gLEYEUgw
l6Hhv5QkLqY+Jf57iSBrzoFGr1/VwhFEXtTvjsJ60R3jM4sdgPbIuaEFfFk3gcKiwmwGLpAp57Yo
i420x0nqP4WKRf7eLlD/yWnqjeJIufURXhKIiA7JL3qWrBkWRXTKQbfhc5YmN5iTpRxX25n3EjvA
lzXkyyTK7jbT7PgiC/9onMFqbXZMjePQp0u9e53ACN6ZjeOheLmiyfo9RJjPAGX35uitppoMLSCK
RukTsFwdrPaFkF1OQMFqmfC0SMXB/iM+oxFE0mH+7SjEvcin+e0ULpdsW5ubeV3nWXxO2VseF3pK
/ddQk6QtHjL0v7Te0e5V+fVSuJaDh9GmYVTeK9QcQ6IK7fOGsrNm5xJD4TCjeeiBjlVRc+meTuNI
oOtwhnmiVjRakE9DG79gDafS1PUhgyxLF5nxMmzga1461KKlE51opALzVuCGXac2DI8+W4kPsk2w
lG0PNY+rW2ZYUpitZFHxeVSqPFWOMdysmcqB8JuYPI8dWuTNvYC6c5nt0BZMtu6fm6UwSv3B5f0g
ioIWElCjrd8z9dIGJa6Or+WbDzs3HAEXFKk7FS5sdsdUwh2n6nZkOkmNS0JH3e6tYwR0qYJ8Rioo
dM72K8bEOrCb94QO3MUvLNaZ2jeSI7ScCz2FMmuF2QOPnr14Sx0NG4qQPLWrbw7WQHL/vqMLY7Bz
R+LHfCe+h8i2bSIH+2SyaW5WbmD/HG54d4QzJQLwXF4ecDfiszs7eQ2qYie4dtpp9gEWn4pl/pEZ
Y1whJh/0C0DgcXev021TF7/s1r3Vt82rksDlTA2vacyUQod4tLYgh9faYyiiYxLSqHiN06fBeG+d
22UrX4J36n8cYxgWl/YiwcKaxkSH0Pud742iQGjvYanLymaCD+SNrw3jrg7R1+7zV/2BMYJt+CSx
Uv1gElIBIzyG4XhJkbU4zR1tPayxN2JtDkf77hUHb9KrFY9DMF6w+BoYjGSNF/48JjBzT8dlQ3BI
rBuDSCTh0kRfXU4JizGOxHwQZzSQ1F3b+Fo/tCoT7HZ2kWQ1VNK1Sd7h22MUiNK+lanQanLLo8Sf
OnS6rhCa6NCP4OhbVfZqM4RPasUsEwOGhRsWxjKDCbKYn3w52Lrb8qH2E5qlewsLFRoktyuuz/P5
80l3VwGYN6dBzinRQ/v+Harzg/jmaWUr31T4IFjfBlfUfOjcfRljlnzZdvMjlfPQTLxW7Y9i3hCL
DGG7hQqTIHlGrWZi1UicFQYhpId/qjiEngYiSIrUhGThbrEKVSF7sIqgL5SMEw05+dgrm/O3oPW9
JsNJGpNbvFuL/QZSfF7QeXiBVeQsTX/9y0brSY6rh1eTeO4g212pM9X6kSMFg7nYVa1Q0P1iqkp5
w/1ECjEyffcrYbj9t9KbG0N5W2Q1InRFUPKNsYTKGRZOOOaJwvStim/AsUxPNjgsN4EvyOZ+0kZ8
FXEdR5m0VE7YbmXbonD9Btp8ASaTreU83nqrzCPfS7VwzYwx2RFSvYr883IDEsIyf+x/sxbdcb/c
9K+FjE2XDwJvUyULQxOkel5J3iO9KquXOMMvMmm/fqlP4GUt3ggIXJyn4TeMwvXGIh9/v/ZPzfoa
muX08rCmCvqHtZG3fthFOSkasm3ogp+a+f9lIFgaqRGxDFQs7jKG4GZt5Oy9NYPVsYi1TVIpJOuj
BOpJghhJtFSaY3EjSNF6bHqcUz2oY0s/5pZ/jA84gHFf29YYCGTVwGdxr5rw3ZTnLTUJVs6JYm+F
0Zqzpy0fprMVbWVNFMk263ON7lqYwpSg+hkymBrAPlzVegVFFlG3lVFvVOQK54nE44lnZGJQCW6r
9Sa2Q1BHXnlxRjI+anRk866VCIEuQN1UZ4WDP2lgY1h/I4JFFjDxwWil0eugZ9bMRxj1KCLfaaZ7
AZmr/tMfufFadYPgnth1biF6UsjX+pt6BTlfRS0X5F/rfaZtP4wZ0PnUWd26Bh8Ysxr/YzTgjtcW
87qeek+6MfjW2Wf0gxmIRzigu5fwoflaX/6OU1uA4vDG1Rn7s4CMUmeZthGBdyB+UIUg70qUTcue
DHxM6DQNgBwbzyT6Eyh51bNIyojcmTwessFGuqNI95I3G5Y2/TQ4j3b8Jz8L033/zQ793RISRT6l
s9M4uRZOVQR7UMD4DaILM/FDMVCa602A3WXMDEbqrtA9xZxFD74l7CnOBZjET+UeLPXmRgAzovFF
CfJZsQKVSiSiCqmAMByuek3rnItwxhQq6AzP1OkUQrRl43NuQ/e0pG4H6adbXnUzjhTBY7HEnWg2
YEVYtps5IfWx3Fwm8xOAAC6JqMS4Rb0bA0XDJZtQBLDaQSP2zPCufDs0Yd1jceCFKeOTwvc2RtCY
itHjC9Dvk1PHPe55L1PjD5SBVPV4FtcP5d3YInAMw2MM//Livb/hmrnl5aexBEH13r+IwlRAGXcS
p5hcvJWYh0oV+wCDQwHKVntmFFNNepHKQt9XcZ+B70j0V4wBaDh6clcV2GbPAhvPshdFC7nesCua
Hf7rRTvK72MGNLHH9Mu5Lmbyu8WQ8dpSMK9VrwkhD60kJm8BRtYhwPdqc3dqdQ/zoQeOUIqVOulj
4GiCO9aop+1v+M0XleWozqcecTdfzyQfr3n8TC4y+G3d+lb10fNDCJqpPrQGIVFw+BE8B6nPv5Vk
iya1HWMuJrR6Hhf8grhlsuNtxhnwq3e7uWVmA48he+hjrdoaDBBYszWkUyLt3veTq9j9F0gWE/Oj
Gd0bgOYOZraI3xmwUBCVPqhBBL7NClLr4wvtTWD80JhFGR4aSGqgmy9gmOWFELoqe0ntpec/A4AR
Lk7JIkH1dRGg/FdZs7JKkrdY36NIFcsWAOCfWR84nbfDAlAijYZ9GSNKvxYMt8fGO/xvSMM3a6fG
sQvwY5jSl0kOoNvVR6k2W01nG409a2n3+qxVGYSl1ZrFPutNV0Z8QtJkcFKW1mJwI/KX+IH5vSHt
hkDBL6KYdG9jE8qQYtrzRUkewtlQHSZK+nVUG2D6qEtNmt6g0dUgs8uL5vkz5YNxJaUO+iVVub0e
YgPR3kHovEUsdEbwXyBPRQVXd1M/bURKZLWIVX43KYWzY2SZnaIVqYpwI8ilFnGfJiAkhNxGPT65
O/Q/xQY5FTXixg8/yaHuUFa6/T0k18ouSuISvmRgx7FuvZjZbyIxhKPtqjtJt8hVy0d3cY5bzHEY
9X75ba7aw1T0FLqfsSjSBCaWtjqrR6RThgf3Qi1H687C0xysdSr/Bs6jpZBtUtqSWOZblhx52biz
AGBwDlG1s6jAcPjAWwMwyMFTNBLujtMASS7yG59FaGWjbF8hXGk+q+9uiUlijTKDkn2KAreeKU8I
fg9KskwMVMylB4rwPcABa9Zmj0Tt8AFUjiEskOP2Bg3VFCwMuwBfu8Iz0+0ylDk4NRMSBwUbsJOs
Bf/PmL5DYCaccKwWHZ30ZurvtORyZ7TuAXmjGch/vkFHK+Ah+oTW8/7i0UOgsdLhtNHyN9ZAVaVD
DQNwGI1Tl4Ff9hCbWJAykLl8G1mPOjVRVFv2QUl1cx4ptYHMECEGAuxxyWUvAqoTker/QSLgeHza
bGGd/KxrtlL+v7k5twtvb/kEfnSdrjaSTIvERZyHgDRTTg+gO+75yuQDWp/8BF6hpXMJsF9Wie0v
yxy9xO4y3EawXICIby200YtN/Fde1sYRUzO5Ebvwb4jkVeOGwUq1LdrKr31KcNdCZ7/uHcAKsSmT
9pP9OS1N1zZ+eHQPRr0ST5eCA12AB/hy7S59v6P0izaFgzw7j1caDEoAsRybOT0VAF6egwVPuVDa
NMhXnDzUph2q18+8Q/wpzm1mU/E/POhrUOJs6dfYIwdco07eprqrilma6Yxdh0iH115ddPKHdjJg
QxYLljb6vecswaAhS3qJaQtwnFGd6o+vCK7tfWhaO+wrGAZyZZ9e2vCLcgczuPUkruDoh+ZBK2Oc
S7ZH829tPDc5Xl/Ac3FfkreziVxRkAIKgOtYAypgi7iT38adqoS2uqxEMZgrTULxUNKcMEnQ/Ud5
dDOeK8fMFFg/KWfaxTpAFYmMsa/4TLihYJQfG2JYobrGBpd2QahHrn4dMVWAQbZkdXWpzKpji013
9aaF2sYgZwOaHoJ6nhfDE2FPdcqHxcAkJFXgckfV6y/1Yy9XY6Fk+Dx/UKBo/aoMPOl+Wj9oWofK
E94ju63WjR4v77d8u0cJ7wKDRDTHiS12FtCXUFtf+oX0F4XcBXREobLP+Kssknr/nOfGHWg585MS
MBNkQrRVUkekEQvvqoX9sOaYDQm5HTDxBXLCQ+9vzxX4TeWOf2avN7rFCATiOvxpSEQc2iBAKjKk
9BsgHwFMMXaxndO4U5hY9pIaffNfuuL/0sSmFcSczKZTNDyoYQ4j+A7yT/amvC2IKHbK3Ig3n5DK
UoCnqvX/aDMWVI7RunSUf4YB2Hu6ULDKj2nZTFN7zIVnTFPP4x5GW1LmWinwCJ0AJsXD5ANb015v
xJqSercV2VBGjK0gu8iBgFVWPMBEcHT40WBSXKX4YTW2FLxlQAJEVpYBIkgMutKltsDOQ8gPescr
DIR5CWJPLJlHPclVKlYeLKE4RIqIRqhF0px/sXM0XAgxdVFKz7NBYIpfdjPe9OsCfuHELdMS3vTb
vQ4OX8DsC9/avjgk+zlEOdHFFz+USlM6chvpE3in8FQeTiw8ygaA3bDy9wTDXtGDO23M6fOBWMcT
apWHGzdwjZh4Wa8Yr0mrXVYMSRAq0hP0aYCksfgEMOrGk1/O7Xb+uuItwWTIRyRfnWcHfwkF8SP6
QCgF5bPoGBMYME6Mr6GXK/7TMwth4PlXLXcNcXs6XsBvL6mABjkiXHfi4AGGffPwXPFABv8ixVks
z3tfyjkMi599FOoGSqvGp5fPxwPFP+LQC+jsgLhES+7/1DOqeOVscd3QC5O+YJs8uk/Jul8curTw
v7IATPCpxAZ8dhplBSUfvoFRoFW1n1fmKniCf93hvGsdKUs+7oLPiP+tXWU01RWe705yAVvN3Rle
AjdUMomF7z1Df29RiYv+gNpVtfjTsC8iuEfSG5coyZ7AW21BDNTDiELDnZen1ea1ibAA+9FYRQBC
aCllT+/jH/9RH9omlS/0uBU6jhz8Q/CbkL37HjItWCk7HekB6jL5q/4F2AQODnIdOWD76chmS9uZ
wR0VL3GWeUiVG2EnK16fRCAXIwfeM5BTj1lkuqS4uBV9pu9c/2xw5Aico0+HuPwqDgxQuC04UwfO
NtEXdp83cShxUp82DDwqauMAh8fEv63xtzgwbgwuSGfojEeMbn1Sfl8S/kWiyuVoG+BI5mL/qD2c
tzk6dKLT8KRHTsibAw775VDb9H4FlqgM+p93s1DhOHUN4pFqc4r6ubOv7k4xcRAmgN9BxW7xwlja
ADa6251W7lIAvPBa/1RDTqsur6kF0Npdu0GB7oz0aDyBu0f6yEcqHiwpVnBjmDyzzpv+k/Tv5dhF
Y4y2KfsGSNa7z4fj9rQN6SnUu8Rj4dt4yo4TevKy2lIV8KVgGGpYq0Po5e6SFg90kz8RCPx2G8/4
kQLPBnJbcCyPubyo9bSHfGsr1DDjSIdrHJR1Dfy2xjdOmwJXHCu5A7wzrJ8t6+Zcw0AwK9FfCE8A
bQs7L40u9qu1DrGZwoCuQ9vi8zfv1xfVxJX326++4g8duM5g7a3zNSPOhfirWqEl1NolaeHEp1hX
nb0KFsVknMRQPvUIPP5Bcv0gMpGp+ZoIGWhVKni1ylPR+LTQmv9Y3f7Lj2GBW+nBJUGyq+RjupGJ
Z07x5jxpkrycrCHCxJxCikRk6XUXcT0c6bavQBmC6uC2yL/WBB8iRU7CdTKXOJ8FvKcWQzkB92r5
mmrqa33qbVqmuLOhUJ7eAuYRb4CY3o1KH1JmwyKv4kOuY3HgMvueQQSD3sOLjM9rOJ7rZaDvEvSI
Rkir0niZmfIUH3yWtaMdhq+WyqKFnUlJbuKkLif6F+jbUrusZg8kY/zJZLhNfzP2pmWURak4c0pT
xuOahGi56WXhzwwJXCow8OJerF2Fxngza1DUzR+Di4DfBgO2jJPeDzouMwAOAGI7XWfDwZbahyZ1
CQsrhBV5H+weWvz0JlL/QdNCFJ/m3E4lOoZKBkORyFtiAsdA4FBf3plyLvNvirvAKwIMLFFGUthR
MsjK9Bjr6X05zVaJ4vYK8h0kG7WJCSoivtzkwqST3hwFoDMUkD/dCQScr9GBEf2d1EvpB7M972Tk
Rv+lCHltN7fqlzru8FBsXeqCWIQb3JOz7LPqRGDsv5C89c1G8CWhjY0/GTx9guhV5PJzT9K/WyAi
tcY+c4nqvSfACTg2i6oUjE567sJfVelEr0PhLx2d6iGjjd8JRdj+EyIPjlhgWb2YxF356kkXIiwz
c1TqaeoruM9GnzuwQbdzHT9Xotvns9Ny2t6ynLRc16REGetQOpMzQ40OFV5dOgE5aRninaWPlyZw
mS3e4r66/cOYMqQrgbFt3zy09Zx2HHZoX/Xfahy+oO4WS+y3+XtHtICtBquNUAchxdM+lt6ty1CK
to+DZzY8T96Byk7n3XIRZuz6/6DxatybDRMSOBY2m4sHGQp20f3Uc7SnDzbV7k9xaZTv17SO5+y6
q9xV7eo8ooc9AJtrCpC/MtahIO8vK3OrV8XJjzjgV++xK/2uTMC5fzifbVvih3pUQjmsdcbfDsAS
7jrSRVQJhrb33Z3HTF/OUNO6Mb2RgKCosx8FDYFOnnlwhDi51dlRoUz4UDBYzJGRor+pceoA+JCc
dyQZYVC8eVKZ6H6OpNfUOT3gQ+J9bDTAn77fJQHobWqFDHLsiuFf1SR4+wCn6bMSwKhk6MsOvbs8
+ggS1Zb4Gt8+7gHN98M+sb9LxPUa263e9lNLrdNHaygUZE9eOMRvjsZ4bvTv1/n+E7ZL+S2xuPaG
MkLicPljM6uhHDjxL+mVNEfb4kTimmYGXWgzu9aLrhFQ4lG3tsMta61gcIpWwFvQ7S1/Ybw0R7dS
Ec0BrEtvwXyMkffp0v0IcdAxMDeL64VZ4nbOAeAjWXPmFtd9WM5siaMkjBRo248ogwIdDOnqiDYD
4yjzN1wWoou/Ea0x6Ds9+U2QxXVWI7IrGxeCy5YdM9dkBMvem51VGZ0MGZtZPcMQFM6pMbitMvBk
fGn+rAdGHPd3GFlQC6xAgtvPdGAP9jH8O7u9W5YTKjEHKKrVYraI55T9mO5safib6fcbFNYAk1jt
wandA9coBzi8Ox1LqSm0t+T2nMHV1OZboYrVqFcZeDyVVHzQkAR7lliKVucxj5ROcdljwKzleuSv
uMqHuUhlKZsltnluN7Gq+WgB4nAHlfFyE1JLtoc65y/n0tVy/TG2rI9xOsmHUFiBdV089S02XkwN
gLGZagkgza/yuVAPTuLMdgZHiTJDgiVz4FKbr/AFu3ZhRBOm8xSv1NqQDOwJKG6ZFxfVc2i1fNEB
HVRrH+Zc9fZiTHt9H5sh8lnhPB6ddx/IYd9Tep22wxApN76kSFkZ33091IpEOYwms7kQnsxuvwuX
FbLiBH9eU5sC/3ZduZtLhHGTd5HgaZalJZbIc1uNU/TLn8TiiGx5EyI0NrSg9jTBI/QZLveuURYD
4VlKqPpLFakAOcPAqKJCBVyoyhXHCGyEg49AaNZ2hkdAT8j5owMFmT7DC6XLso4pqKfn3eqWbB7Q
VRfroRDYGkMOd6PMDmN4k82cWmZRZUHMjSFG16nBZAv31lG6NStGwDJ/OP0CNTUPDVG9CU29FMYK
tA3cmAY2KkldRKLAv8cIsagxtaOnIYAsaG9uUanwSvDi/5TnyGiIZbDSyvefESbMgNnb6CRyBcHW
cFqvv5iKzsraeRsMG2nGox/AhWoXU9Gk595/jzKOmTaDZ4SVFIcPqDX0uQZvuG+yll1TltrHnopa
nVcUvatpiwZXgnXtc8keQnzJjMgjU0aAUquf5/fPVXZcOPFXL1D/ZdJYRvPQ3VdH6/r5FCKUDpvd
jMPGhgwer15d2JFvO8vgwDFnfqbO/wV7WciICUz5rBJIr5BsP46fMnGgS6/W/kFXnOwDceUhSsqz
rp9IICMjOP7CW3DUdal+DmNV1wMvrGYQbHdMOTpVoDaBCdO3rMUPhqbchrj0+iMuhyh/O4Q5kuQt
kNoKjwnrC1fV8k1Cqi/pfR2OZJ3YyYLC3SRT3SoSzC88hCWMsZ3MQg2FKIuFkn/kB6SIxArkJ2el
irbmh6z+klrgZstlRppAQCRzVIClLxu/sxjzwX3qmVP5xhDUBQ3ys+PzLr07vqlcBcefcind8/As
TyWqRy+iVu+WzExPW+CSgZFUosYfvRp28YSqm8x3paNMYWM+Nfy8Wmf5hDu+pKn65/2M+r7n/CLT
A+fv2axZgHC6rAHKgx4jdAwcwc8fNhOHRrZe6gqQGcascDUPMIHE9OMCMbn7xBQe1R+deYdiUxYA
hRsiEKbxMWyObEt9BC52w5co5DqaOVZMozygjxX0vK8tDneF/ATvs0GxzquGs7Arjkh3IUD6FySH
mFKQt6Hk7mj1UrygKAdSNHOcYjUe+xRaf8AyrUTfaQONTRSZ1h5gKQzjRCChNELrvs9goWDbP/ZR
Zy2rjXCSvAIBMj815xSDHOv7d6bod+2/orrrD1+vqyRwD0EFrzaQ5x0BEqO3vPM67lEhhRXkrCwn
+/5W8JCR/NAsiHHHJpZ9V2Bbccg2K/AYFSLYUOE/nRM5C58ygljlydH7q0g1nkPXapTVGVi15W4f
tleN7GgbJCWOWGlj/AGQQAyF8N26/GoSjGuP9lU6ChtpC3monziEuUg0auSMoR74u4YRRhC8Efkc
MRhmdMyMmNFkq8IyJbT0SZFrMJQyjlbtKG9ajj03LYq4qxTnrHGOqYgbsuwRXW5XjIIYCxM5z9fz
7F5Bm5hU5v85f9/8G3thI4KISH8ZYLf62wM45NqB5q7WLd1ZKnj6MX+RxZYzO5nJdKX8BeFk30Qk
fhSxGJ1CxUNMG49dVx6LnaF0QpQaJ89z9rzFNWkMqQ4N9ZwWX+8Ci1E2mXfYPX+eQnzzRrXOMxwo
WJZR9/GllH65pEsdBRfJarQbT3vMt0UZUCd20kexqObdmNS+gHRkGC7C36KdDjenlVLm/GW0rYJT
vBPseja1kFjHFnMbcxdcekORRdQMkC0z4UnIyQBlMBvcE6PhB1Kf0mK897nNQNSwDwZPulDOkOKn
qTxSDAoMAKvu2qiCYyNU/rBOAWLTKV+SIltqa9YGbYCc2WSpgc+WWUOa69qbJevMrA0ivdRs/Fut
uDuGhZxWlqipu5k15fPhQ5CxQgm4Tsvz8S5ohD51pf97cQv8qC7psXTNTaSeeExSLKWsH9UBZGfd
VAhtcZJ9bGmwErZ6fLM1AMMYLz3BkUWnuIiQMch8XgA27oArfaVRdDV71odHKkiv/cPTCbA1+CUE
eeSK5xqcuTQ1IUS98D/qiKeDSi1ZtF1jWp1UwAh9VNxnDIeY8kEefOrbfJK6spSt8RUjkmAfD2cl
Iw5736A8UzzKAKJo4MuQVZSfrBMy9zpDB0bhuYLdE36F24lNHTpNabEtNYb0wcwPPZ578xZ74gX6
AGIY931EpWKsSNvwGsfJNroVdA7IxLBeciJOZAlJY0Z/eA0nryuMLKjCR0jEuZ5761k/r1yVccsS
l+d3V+5IqjSK11M0reRd9/LaXE4DLP5BEQEai9aB+WQB+fw5AGTeCVuWfzwKAFskR8pg0H7i4140
64CxRWJ1t1W4eYHz1Nu5eiHxmSsNfn0V0pCV5Lri0AHAW8BKAcphv3BzVtnrMxsSAModrVYKJ9fG
vIc/h54/rGFcvzbpgJBZB7PU82jeEu66oHCs0TB1Qy01dwsy2AQRhL38p3bbE1GTnenZ0KeOpKhW
eNotlshZA5oyiCh4GSaZlldOYbZP0bizZ93yuLDnhv2T63RhhOjBHXRigsfAAoBV5anYG7bFtYzM
TIiDAlP7gsArb/jnINppp+ip/zEtDZRSUXoc+227PBruPEMt05XUnl86RF1b7xz+x00cPAa/Rr13
iabwU6VLLmXn6bkdmvGKk0yZHeyrGPRt238fc1V8n7B5761qF3gQQNUNz6Z1KashWOJM/LQejVmM
vzeqUJAshpDhKQczO2mpJWYY0fkucJ4UO3MQfYQqpDxK6s9NVqZ2/op8OAxwCyQU/uSnnJuD+9FG
WtQs1GMgmO0y947zli/FgKnRkCizMKu0L2/L7LPvJ4m61rDCKD+qvhj+KXkdzSwIftvRpNG6B7Um
NKtHH00x5WjoAtVhmyTczAH/xRXmjHIDt1vi3IKO6wzLGXq8eSpEy5ZtbH3lZ25oKaCol5OvyfIW
Hqpv84ms2PmsJfGbydh8V2hI7EY98thEvx91ibGMZixPGBJz/VuXUP7GGnHMGLRCH0Mg5F66aqF8
jnW4uoKNCD64ZSJqwAkFbKb92JMxz8eS/hxDzzixLbJlocKhXluKp9ZJNwHizvq+uz/d9oyVKy6W
UVYsthxxJC3VtSvnx7cAtFN4IQj3otdDWnWCfgohFivys80zGkwtRIHvZ4d2AxNxgiTWPVsXnDtp
utSpjXc8dw+c4yekxQ4k/seapZrT/9lhtdbbBE+RssyrP3/cIv8FWi/uzD0ooW1Qn2pzK2Ksj/Vr
5RKBtEJo5U0/fJLYf3uRzEZU2yjReWUzTBCjM1a2aCwX2j30BzyxEAj0uvhTss8rLGpn1wBVumqv
L0XVw7BbOUye4nKyQbyOR9eJhzIfsF0N4OKk9YJau3kHeptxAcMxyWiRp/U3cKF8Q1Ed8cEpSPD9
1S+rYKsCnCbJlstNZJ9cQNygjEJPOPSVG91hmil6BxLK5nXLwxxd/rn+C0Ug+V4bBAbB/Ocyfl+O
eNPmN5XnJ+p+AeP8EzBYUXJfQwcbKlk3nolbmnZt1TYTtaisaBs1DVUx+CcQLgYgNflcsNKWfqRt
5DCqvxqwuBhqKVcJtq9ioZxU4WlziUYp3XSjgjzSEc0td9Eu1NaG/CEPherfMpfAGDcRW078pE/Q
uRKLqfTXzjb0xeopn20KaHxgIMg0FeP5CFIVREJGHJRGFNPjewOfQkLz5MqDLjJOrgUYzzMeFGP4
aWI9F/8el1e00kiOhNxJRDrD0SyyI/ZzxuZ8IUx3FNJPG518TkycW8oszLYX4WYorGbUt9QX2TNe
rkf3aNRqvLWqJVUN662jExJ7+F2fyGPlAN7IYuTQyTk5eYlsk68axHSL6jSP0YXrATQlgkZJvW1J
uZVHbcq5Z1xIO3smP3JIPJDqxJIW0aUhqzU0KmrnuBhDg7TQzAUWSAIDIr2dQKKEvJCym8tXbS3u
iuMNsMSoiS9sDBZYboZ7AmfwNmFkMGlrxgyN/PbDkD1IWCvzkvozmltCVxTSdu3Zxgj6vdf6hftj
tpVChuolNVZ92dukk0XR7t7R6+igbt4gOrsbDWoXLx7jOoOd9DJxlwn8pCn+t7wCePiPEoPhKeSs
BNQBmsNGcWgK0IFTe8I1WL6O8Q9OiJd5p+dgtu65pKVRBtERWLLzobM1AkNYDOAQqGPIS35yGn5t
ykGRUA2PQ2ghUEUvhFl0aKhs1EHerhzp4+d11zxFtiD9QXVZIU52p1eyfpdIDsZYQs91VUk5YunA
tt4BiMcXbwTgyPaV/z1zx+g3zeZ+vYtUrz9MrcxTNI4ejM5UM0UEQWnml9hmtLt0iUMTjQtGytrD
590dEajAENajFZXlRD1cDejeHaqpjVDXZNBODCj4DzveyniX5XZIfLXqK5GhKgoCzdgrNQOm9T+o
LMp3O8CCxmUY6am2vjYSWXDyUjCIrD87icG9ybvIyIWaAERALNpagzM3sXwne7qg/vlAPuYJCFpr
Qez27TC+RcF9d36/WmC0QmjS6d/PC40IdrFrhAWMSgl8AnwdLzEdVbWmtMo60UYy/cA4eS59egWg
+V/A7pIVAOPWccQdhOT1c9tjYH9K7DpHEK/pKC9izdYSTa/Ipvl0UTE7/LhN5fbfxbBFsBHP2+fB
hQ379md8wRGZUE3oLVR9HcV9Kyc956TnC7AM06hkbDRwmFXKcE9cFxd2V8xmazVy8FApOXQgMm/d
WpBY/ss1vwHiKuyVfEIVeJPekrTui8y2Sm85+ozNq2DK7sgqXXVhpVPjVglp+aSaRhuwNrgANXwq
f+AB9f01ShO9vQ3bJnXCX2qMd16T2foc1DbmnuJCjrvojTa34kHdx4+Uc5SR91MrkBaxHgW++FPs
gBNSjSiihAK7rEtvEXs2CvC7eOVKeMsKDcbo2Uv3RranIYGv2tdU2ssmcfRd7q97bQ0hN5wiSba3
DULQtZLISbHV+S1/odh7J/XDRgR3HIlzNlCq7chdlwqaf2em+J3WocADI+fy/rq2YEAc34kuftST
KxFI4vKMDM4aJvHj1KvJug9pHLw7m3a++nXz3/QQhMhJChMYC0eODjmZ8oVQi2KzXacyPHslPqRU
bqbMkScujHfU61p94kN4KjnWE0MszTw0uQ9MOmzRRsUVkS4QofyO7hQKn33QCw1htpwxd0UM0zHq
uGCRTaL5F7pvO4vj9DdT0ym9tgfkFP3Gc5XeRkyZbNo6NgOmV5gP7K8sSVsUf427ft8f7ijBZiqV
mjnrv/OIblnP8BIE0tUqRt05A4Xk7cREnDQpOIJUw5nhnULQhfSXvTmw4wKwn+1lwjvbBqpUodAo
/su7kOTRCsnB1g3k1t/Zx2uoIaDgRLfTjK+IZQasNvB5Rc8uGoKM9cbbVEC/SCyrQrPYLlUXZIkZ
Cis7NMpFmilRpTvSuuy6ZROEFhd5rJ2NEXK7P1j93GdjGOMC5iniyhI5ppqphhSr1kCrj/Nr2lXS
HJU4CTXmjjL4Kd1TqPwY9jmPVDuTgb2utZ9vwMCPFT8lOOAKW04O1lA8miBdrrBpMRoGbS0BvdiY
UvkuZJktplDonDw6s/YsMGs3VBwAzEdJOM5b7fFnTM7QCdbch9A/VqaQD4LN4qswnhbDhzjuSp35
XheHWveTW+aejoeaaMNj50kbgNLQsTOVEEN/zEXLvJ3B5iP1Auzphif1zbvVlbUnkKkBPOD20164
WO0tiPadz+Lve/zx6HJAIwwiFkbi+5nftGGk7zlMa8TffAA6o71E/ZsJr7dJeRER6HesaougVOv7
HpPMTyppXgyiBKqnBv5dMCo/WSAnBEC9glaNdbd6dcm3bNQc2agId7iI1vbnIUpo5IoQ3pXwO29Q
uCyR7/sBo3mLQiRc3CpwAd2rAWMYI/8KvghfmJMmSUQiPXgjoSeNOuvIvU5kU2zhpeYoW0/2+r5W
c/OigC5Yfwekh05i7lk4WC7voWQhTH7eUp8hK0Lbp++JtsxeTAav4pk/0gKh4PtBn38sY910rSgf
fZ2trrfyhN6i3zOtIMHXyoMpMial8XzyAhMk8NDQFl3J7fYVGW54HppQMKnCDVWIBz+wV6qQHfJw
Vh0mOTq2wjwNwPxGHnQwXyZpsfXRRna3e5rVsxUuTvsTLX7CRB2qtReuT0McrCNYfDnVwonkJ+FQ
suPC8StJZ0YjpICYaGmuqHw8fs9uFrX+fzXANi9Fr8nRLnuhmhynhH8gXj0Q8788HajhxEXDGL62
ZUBCgfdxNuLaOMmF7UO2vZj3Ohk6s6iowZbQB9YBX6wzcpnAxmhtvsAv/hQGXAj8gLekfVEbta8n
sreBzu4wBYBN6Djk9yXR/DFAZL2nV0QmruaE06tIzuPsmAqYy/o4h5yZKs4XRejpMhkNUrrKeBC8
ypxAr0YJjcTXXdDfkuuY8SeeOkSXg3B4bBhBvMGtN/pDATjdecs6SbZoeFo6UbFCsvgWp9WdCJAd
B1bwhdNGTWkR5QZUpoEA8FZIrc3U0b4vz8YhiEqc5PDwvGlY4OgOGREb4mx22kuUKHAEefXiNyOE
lpWz791U/cJS3ysRoWwwLPUaeiCONJoZxRwqh8iu0iztKH4rCj5MmBo7eM9ygOl9U0TUa/VvX20O
8RT5gN4ScZj4IpVoXfEe/dTwW+z3KTnUS4+xy8bLWP+D4CWUoLY5VAXP1/f3jMZNnvJ8wV09JaKv
xx8CP8Yh0EKhv/NJadXt3K8TelNgV7qz8Rkw0/MPbimvKSGFtIIHILXKsOjuWGVcb27POxWsElaQ
RBCmIxKthTmtPBGXh8yM9ASuZ9dP3S6LfJjhHwyqTRFvHtY+7MPmuQP4njtjHundjVZVLSsH8UpA
M/focw7kSKuXsKamRw+xzzhlFloVsdClcllocnP8EhBY00l6YXJjl8qRfFd65RSqe3f4/XsHs2oQ
8eMIbD9Dw6+W24ZyWPbL+UdIm4aGeUplZUYUVXEASa1IOzmJmj2VL6OM1sy3Z50I/CEZfO9AFYFs
njIs3cZhZTJqk9dF8O+fZaxOnme8q8c0pD6i5YkAvL5/4/0S5pJlJ1MNPtDc7t+8wcVlA8jVzTrm
R5Zl2Dh6g82zRQExPvqR7nZD5ca0KMAwgelpezJQybU8dj7r0pQ4Y5Nkpq2oEWtcAVxZ01dBDJtg
fMqIMqRI8LW6AhJqBGdOSODZemHYw6tqaXQHJgqiQa598bmL9Kd4w/JBOzz6zZ3lastZWRIiszVb
0EGQxFxB9vLVI9vMFEeuUG2doeumHhI1NvnIG3LPbLAtroCfJyoZv3ZyQmvg+jOl9uSi9NSl+ndn
5ClK1r5upEdOT9mr6hPPTb5ANV6aw4S0S52sdudmWlvlw4FQyhWx7rVDmqGKb9vrL92r4gs0SuqC
RWZ/dhU70TYiNfVhVCTJIGvr+D5tI1ybjf2FtB9hDftY5SAof3TDwu+/IGRT6E53dmfFbJ4EL/7d
MuWdlYuaJq7UUaY2E7oBMhi4soj3W6UXE+lPk0jQzhEMi4C4xuR2u1c4XDlCb7o4Zl6iicUaWB+6
0UaLxjWV0XOQTd8bJ0m803Zo16EtG9TK6hjt9vClOntmLyyOmf1eRHiy5Cv81Xh57nYavlXpc1Zy
wu2i3O4WzNfTGjMIaz6XG6FSxuIY5orgUj8OHJgMcujoL1yLeUMgmac/Io4gqHGLR2ej435IgGB+
cUtOY+73a2+5xHEQGhhmvoGAUiVKvj8TiMOO+zH43JMtqdFEglouCMq5HqA+udZ3HnpIpeuKXjha
V4hbaNvupjIxqr9B0W5l7Gj5b6FS1THfSO53BPjlECufxSxHIPpyoqdOhhOanXkq2dKmS8LUNrlA
1BBpRa2CSEqEgawfj93MxZA35h+YuO3mxm2FPy4WhRkuAf6MkaFmMzQhPlvcsM0VgODIDxT+9E7q
6Eh3bvXVpUdFVirbKDcLQHh84Ij9YtgUG02OMvysUx/6TYaGsepmL4uwPCv1zCtv6/cp+N1rPUkG
ipZIQgBFtWjdjKeVwUBMasEP1ZRLV+ZCkOLKT0hncHpvtEX0v04SSNTmubKqH84gWU/fvsPEtXZR
46+g/tbgEnY3V6I7CQS1aR1nwolSaY/V2pfr9pQL1bIU+tFVHZ4OQv/bkrA7tqlcJ2vvlUEQGiOH
djQSc573JQlcKVyICvtWQAmcB2nyKyBgzB7jBnMEeuNpyRGJa0w6Bwh0oXoNhfrVl+Tc5Axu+aQs
EEpdze6eOCgPDkNdFLpsyPnXFr1BUFnGnhxwa+cC3wExjW93qiOPOeVgVDNn73v9dxZwlr4HaXMX
R/151MdStuZa7/kmcdVVrE9EszvyBolL7jt2KjEU+cAHQp+aQqJXAFg04fiPu28id7ErFzzyzA6b
4DOb1W90W1/tbZUN2KYt/eWypT3PcXNCY/HA0Ch90+R/xuooxhwy2Q5vJQKjvUWlDJ+/Ns//r2Iy
bCanNlfP1B9hhwWP9f7CNc0gATXWMqb6SZ9iyMTv4uujnvswr6tOgfpHHhHvvUhLo43dSilfo71Z
ETICs3RGKb718lntoZCut87LSuVjv/E5yzaNUhlPPSojoKcpPPF3catQUP8BmG9BwHne9g1TrGdv
OlWRKT3OjfhETd73cBgDSK9S8FhXU8c+JE14BqR3qHGd8iQ/YKz74hhs6d0cDE4G3zgSiLG6zUbL
4riCqiJiMyWlWF4+cQ7SuF1aeLpyeTvKRsQ6XD/mrNJuT/BuOGQlrr/h00m/z7zJ8ux8vgSAImip
l7pdJIKHjQ+0od1cJif0vb9AhkUomgXUqHxez0jzkfO6GKEIpc0NndIpUOZlGpUKfliuyX/A/3AT
t02NeAXtmEVVzC9G8U/GUMuMKB9gnDrvopDndclxaKTqjC6j5xSq8UncDPMhoXuJpnt70CwNZ7VO
pPOEwg26LcQvIxFW1v7W6ymK230slc9n5AfOVuMyhtsFwI9a1DL04el/PUMT5yLm6dTA4CxPvHwY
y3SGDVN0zE5Yq8gz7bsaQtUIj4Zk99564FXBWhNr+ExFL27d0lzyvsNli1v/wy7qrtvoIWTO9Lke
e1WaGQSBspgH/YWUg9SBLZLlm1SkoQh92zYCvS3JCyTHtn0bahxSUGCwSFw0QRVBEOVz2uGBAYO5
KbmHn0aqXWSO5NenO/yoiVORsGwXkskrJuycrtAgHYGcMUFvQLEZg8L05iIdce2FufaVpgAkTyxp
/7wNi6q7oVJAOMpsGJuvdVUr/jwaxMQNm7Yu2Dxl8OaxZksxu51MZolDlJKmFSFvWMiiGWfnZeS7
67xRPpXMeeT1HqKRS/TDYWYLDfMpcGbpI5amWbh92cMxgf9pittoyUoTYD0mEeGYW8PVb+t9E7+8
o5V2NUANohK3BX5x5S3/6nm6TT29RGswEDhKDxN8ww9+2cpjbmS2J4PZut0w4WvQfJu4ZkW2LbJG
P0syX2mjY4EDAkI9C89I9qvy2fDrWvL6ldbKAkFImuEvy602rBYPSUS5qNmNvdU8F7qi2IWIrbUg
Y1017Y5Le/y3ZiUycEFZDRW2JpA9FI9p1kRiASyRcs3KlCt83xnJqaSXY02qzNJbal6FWtjBTqRq
cPSWtflG8D48gGVXqk4KVttTnCucEM4dDtqJVn87dd64MuCyrBdMbryIWmGuUhPDepxvVLXHuRt9
bzh6gP/ywy0achRdMQIDTu/YiunocT8JkSP27GHGvhPGDuCjziiY/z34liETRw1XIkFXLxfZppqu
8MRqR8+oedpEtBuh0HrdJzxkQa4xw4uxPHA4U200i3Lo1cuTNxFtH9562iHFEVbMO4NtRgAxCZDI
hBfp9Eif9UDN6l9dvpvogtWMdMu2bEbemSi9nYJwXLYRsHk7PAHONpBO1op0X1z0OdgLKklmOP20
9Z0+fBplm/1tcng3xea39HwSjus/4D5WZllhJl+hUD2BJaSWQfgkGsgeB703erQ6RSi94/K6VzyM
O0WqzhL1jNrZuM2FSYyb3OVTHKRdxIDRIWWAXRuY4XmCTjBOg65hCo7xvI7K87K0iVP/d9hOUMao
4+ImwjfGEnsDjbkMZ2QpJc6z0DbC3S0ypuZKi0KhdUNSjyjDpSIVMXEM15C3u4GD87HP46Bv8B10
NF/u+BcLjqMzmZLYFArOjWwP6ukxZfzkhyT+bwLMJ85De8XyDu2bRaO3xHFDL5FVWQEKMUKdbISY
L++N9gtgsJ/KohpaJ3SC56eqy3Ka5HDygYG73LmmSkEw/M/GraidDyNhRCs/BorpoLsvRjBJiKJB
uFk8SIdfNq0nED5LfWomOpqrDl6CqaRUoK64x7lKqWBNVQG4PvsFvBruyld6xiL1IV5nXoPiIkUS
uUbVS0H4PsaMm51+AJ5AM45OnGRuyAw/AW6reGGP25NKURRSpvONnimLnT9vLx+zVFi9+i824Mbw
OyVqT72VonnLsq7epnb1iRncDcOb7N17cglrVLKC3Q48NctyTCkGXQbD5ExUMmnZef7dVzmZGb/5
UBs2bcbed6vdx0A1bqHqdnC5+tO9JtTWYpES+ZXPeFm0HWbSDsHT4N28zh4Pkr3T2XLs0DSMs79f
jax0G7DHF6pttSwTLMzM+iQR0JPSkkV2Em89rc8Ts2L72fCOYMkV9i+bmMtqvPUSl6muGlyXBTrg
j/t87YAsZfjipCm/LJU+9J3m+ioqbrcyc6KuddJKkuJYuj6A1JVpUEhXOHDZoxoaVKpUb6L4A6eD
3h9z3SQQOfeHvGfdvnBKLtdTBxFdr49aPsIpC687t8oZPLSLGQcZgtAD2I/4e82d/L+IojY6/Diu
Vx5h0txbE72UiV5vu8g4wP6yE1L1vVgjr3qwz2GUjKaoppWrNvNH9Mvejmaai+a58gqijUfcO/bA
XJtmMl1Ud6hOxJGOw0+2pesyyMTyXtMcNAkvcbX/724oBU9B56hS2l51A2stfxycgJQIGu+Q1ce4
xlHypkohZq13xvfnIKR3X7UTmt4wjsiQV9haiKGhgyagMwGGo9re6mtIDV/U68XMEsJurmMB26XL
mXUivFE7NfyJ3NwddrZBB9GwKYhlHl+Ip6qRpkjtfs2KLDPuqNvsjWnf89LunahwgxQaoIse+F9t
o1H7Q2uccm4KpeetcOdnd21NFtkMs8ayeaGbQ0WQGo6lWpdVopS3TU1Y4XWyRqhORvICqhbL8A/T
MywwjQtM8OAxyksNQuRag5Tg6fYAPQ9/D4Zddu3nHsmmBafhTSkcx126fo/nJWxmfBOCNItgbVJM
3psHR3n3YmuDsTLjYc895o8iB3JEVO+NTokqGeV+Z2g0NhOjJilfVAao4SM297KeAOUjJl8iT/zG
E8DpEoFB+AvIXTU5XRvTmu8+YrEj8xODtkmLPyeiH+2g0qFy5EjHHfJ924l9qfRzzwgtoc8K012k
rSjeDUtwc9+XLiiLRWoiOKwtI8GPAd2LVykSL8dYOYS+2Wcf+PWBRzC2MFMTsbTqWasJ+hYX0Ed2
sSvJl9E8/gLLajtQDzFIuFGtcK2edizei57XUTYbEnDeX+OdwQrLTZ25nPZaIGgpIJJqededuaWl
TWiACM3qt7ZYZINLwPUvH5xbLWf5qknfVqh7Z9ox+CECmapz9X7DQImFHpQ2Q087f1S7H+tQoCbU
MG/sfhY+XG9iERJJxjLBZg5J79/jUjDYxxOpBw8gQXWENE9eME+wWxO3+1b48K7mTBQg2RxpElWz
IgHIWNsJGpn4pUxEQEz6IWiBpZN5kQGbOOtsbOXJ/WI1lRhb0hX8mYwkuzuNejVRPlzvI+SwT8wF
F2ADla+xx25uENY1oxSL/XF1wE9uVK7oxWOUAZhKw2L0mQBhW9WCqyVQGNdFHDRn2UunmlnsE/s9
R5DJcHY6qlt7XCDZ2j/tAS89vCjQoozybYSymkoeWkSF59ItYVIs58HhzK0nIUuOq8QKi3hJcGDZ
TQPUOVzsrqc9f7Jqvq1Kusl3j2au/J4gZJc2r15wn2aHNbCVn5HZ5nv0TaxtTH08gCerRIjOiSVE
lBbCORMlucDzivS2wCYVnQgs9THb4TEGaw+LLDSJo3eMhaRUDTLh0Wu5OyV5ZoGoocWISMZXJ9z4
11AQTjjrYTjJbWydwIY2EFvsN6hijmfzbOCr26vZLLCCFi58bHWX3p16Xp3DjcCz5pcKWc9aHrNK
Tnqp57XsRx87zrRfYEk3/kQbOl5ell8o9AH3wepSs5QanVRwXugr8GPfr91ZR0L40JA3kUnf5bO7
neeyflhKDatheGnvkSpIzoZZUaaPkqELOnyHruK+rvjVuunmT62QVLHvQfKZMURNfB1CDfQvRbqk
V5lQTiX6exzxf0x4w1S5Nh5Z/gBn0gTaFZkTYAb7LSUDA5zdzdndhb3rWnsvHU26nDfxp5LfcARP
uLk0X8yHvaXFERtT13vrIbmFwKHglVWx7W1xjXTPuVFvAgIo/tpBsJOQkelHrPgZyVC8s9kdZi5K
z5kZN/9wkQwzLh/tBR0R3s5W8g3ybOnpEskdhT2bgQN7zhopCO5Wzsp9lciDY+9mHpacn1HIKD1v
dWHY95wmfgn5W1N1y3g5wuGSRFpjFRonMPKiawdfozddXYBseeoNuIjJKqBP3r07mdId5IshTgBH
u59pfgCyF1LFwM7MeU8pGMEpdT2WDKZk8tkiMnEVwx8iaSDOTMfjog5RzgBdc0ogPPOUsV2sErpC
1kPfBjVNZWzvVNeh2oK5cZH+6A95XdJfYPPUtidnvHmH5P4+4ySPCghnmDvTqWnfFvaFlnilGwHE
TSQRPB+ndV8foBlMLd8r4NGYtrCSQJuW7tJJMIY5OO8biIzmmxElMSftdatw7bfzyVoou+KimWym
ipPdA8LkrTG1Z9pLwo95VaPkM8LC8TlL2iUKfKCP0sblVxSwKtNm/w3Xe3032bjmHlIpqr+gXn5r
2c+XCaVxhVRHck6DHpzDLh5IfZBb8GXfDuliyFHGj9Q/BhvvSve96zHrbO44xy9RQOvbhc4eobMx
nd2wGc1/zGHxZVueOgAJn4UqdLaA2DrgYTtZdArC4oa2LTdmPgpRCkMgXz+NV8Ku41aBLzD5MEVm
7dWH56L9nCv94OTwUvP+NNCo169n+klMbZ0B3FyxMFqbFupKt34AlaLX3UFTBrF+ZBYJ1KQIsd5B
2+8ZAJs5dVy6Mg1tMJK13m7FOfEQJut9sambKb+K65GMjKLwH8fp5qRUQA5nUUEzuFimvt6nWt5l
RLhqt63sKHgZci0JSlz1G4xe2jj5CAQNvuKNNbgh+MijvcBo7txFjLM7+0ookMXzAPdyPmnBSm9l
wSe8oXRMu05UALMXtsZVcay5VpQCoY/FC3U2Ci1+Hyb1llexozc7iqk/GB7xeLVzqWvFolkxTJ7f
Zmyo8S9+8qC3GbCvH5FPKHh6j51+iwrJulgkfRVnYgV1aEsW8aQRNMqNJK6DHIYpwwXio6iH5cZE
FnSP2L2hx5k1sgug3vCP2PpJP5v+pe9oWmMDjMa42KGlZxReltnjKpjoUsSgzgILqTlKS7twbr88
qYIcwNeuG72jyM1C0TqzerU2VKWABu6eBLG68rafRnUSgAaTCH7Q1UHEmEem6V5msopyqgerDdZ+
CpdA4WJvIG5ecs5zCxl9eqB/pYdMJ6Dh5fI7D6LkQno9wzYdPGksEbPmnntEB1lhlLcrK/p+/3Tk
hMPDpGxnwyNMaJluqrqpBkM3RUEr1HRo2pKTNsi6Vpr+zngGOCbLIupFIV33UDL/qIQzKjstx8gL
4nNINsiTHncmqPocLyEzZd+udMC2qtMN1TMBIt8affYRm5wlENUl7jsPFrJrzt7G2R1Lxtg3tzaQ
uqtKw9HpMWZCcj1GH8lLrGyRbRJolFJuLPJ2q7hgqmD2dco/AioSJjGH4QSt76H0VnfvYZgZmhh6
aBeh1eOg1MRADqeccLQ+gJ9iT4AtwubXCG8+6oXDVhHJYdKrsPqFFQSzWYetKY08Lm539r93c2rW
lBBcvIw4zxD/s79QvTjorEZ5pIjQSS8V0wS4p0pfxwlA6ANZgR175ntRzikX7mZ884BCP5rcxTVE
4QGURyIz+IPwpW3L0MW3glgM7rD76T0DC+NIlhL7qPoP9zEDhw6ifaaq2qC4mFgKNDJz4tD/8Tsl
nBF4lopI2jMbra3MWjCIQO6POC9IeH5NigPmRpL8vaEpU0kY3ZVyIs579Cz2NN3KsPm6vMcPoYkm
f4hh7e/OngtzLQBEJXL0liT5MxSxT88XJSPxSC4tfZYzLuveDXxzPKT3SZP9i9o8P/9N7NJQjMwm
gpZxlK/An7KABHNg81Zs/m5MGomOBvGn3LySHN8S26uqMUIykDxD1dmXn6lxTlPQ2wecimWg8Kwr
GBhv75uo1MtgvnhYQ4/UXTUgZxzItbC5TQkl5ZBZYptfwgM7cbqz2ch1O5itKtGqkWOfD6n8S4JZ
twiO6bJpGVEGeTZens9aS/hrQ2oRbkcuW1/B+223nJriHZcaTTHGyONN3djdzq11G9XpFW0VrbYE
1tXN4J0Du5wFNPDLeUzuFtQL+Eg04otMeXZuNUa8JjWJoY2JCi1i66eNGOYozuxDOYul+fNTQYh2
qVDsE8aDHktTxv/icuYW/5YtQh0FvdeQyvhS3ROsIam5OzXGxHHXcVacTlGdFjT359YbwImLHuLY
SrXg7GYmOmpSBo7vWnRhcYpWNoahe4P32N43J+0hq6JAnEzsfcMwBZV8GCauO4reW/IcAUOtd7OB
SGS2p4fqmOo47cM2jpuZnJbmfhitYuQTS2h+roZIW62+TsdeXVqdHC0b/Zlyj5j2KV33qoTdvf24
/2c5rw9JNLUKKrywFT0yYiEz1ErwN2hy/Q8oTfhXxXDg6wPCPZbAwZXkLmh5IgCPOlTfnV4238q5
PHelRRwwdxmr/vRGDhBfk/LOymAriRwBkGMt5tmga65k14ITogCXeISLoaw8AG/w1m6YftlJcMDP
khgx3dIfEQghNEgSE/aIaPv34YQmBV63k6O5PMkFu5HFYEK/+Wz/ZnsEUVrtPCywAmnM0eR6AZsc
Bxry8URscSaJAo/WVMMyJW7CshpgvZT3Y04ohTMOKDq4MIA3+o1wr6e92IWT4Z6GlPDkxBQF3dpp
d6AaywRTdQfsBIyYwz/AqVt+6YFx4/0DqooKeV5ShnuTJmlhxqbhYOCDXwWkHKzvdtexBanQyuVK
nY5dqWhcaWxeKbzARKskMZ5pqgf7O6Ey+xV1CMJtUFoWzRwatWnH8t+Ejz7mRLXn9rv71xNWFPCt
XwI/NDaiGwzyMQH3W9oyM+u8ld2LqboPukb6kwwNp/CJpyas3fYYuHgt6nYkb1Mp+UFDO5Yw6lg4
HPIJrnZksGhhQ25MoupyDy0/2QAH5TN1PqmALuzD3y7dtSfm+Nyvy/E+DM0eQSDM8snqV6vJdBYr
3CpxbaN6r1KKZQHL8Pxoydp297IUb2R4QTeZ0fZ5nHCCBIGZ1n1eq20X44y6xKZIK6mZ4m9FQ8la
jGRgNk1KfI3RUhoLxNmchFJCrrqZMrUhX5Ydxn3NsE5q6qYmoO1Pn1iWx3Jsy+jqdL7KgoI5hovY
gm7lHS/8EsmOMQ0BmoYn9ALIaTC406nDl2RXOfj++r0XW/Xl0sa7zUP8PRr5p+Tv/6UcFc44+xfL
M368gUohvcn3bY3ebtjGFJnY4A99ws01kNR0+40LbcUppiy/cgYaDS0L47OlFFjl+vm2DYZOdSWk
LEXqHRxNq+gUBIuNf14B0I4hBpOPjk6by7XHPxQeqi00z3PHCEDyLnAEeSgMMHuwl1nVOWxEswxn
sLAPla4ahlgn5A4W90GKP7NlLNypP7cva9C53BN052YTePgCkmx8dbPps7muGofff1We1AUQ1JS3
mriL+lA4rwuJDY4HVqaGTh4GerHCxNzaSY6r95lPOYRS5gAPfXS9Iq7b07x8+UaQ+wtvuWlMUorS
uabfOC6nYqTa+1uDR+PF+uVKUTwb5+XHgbmQ0RLGRMU1IZF2i5VPF9z3jBP3XLAS9lzRVEM/W6bP
zkPouCpUkndGABnnQN/OgJl604RyBuX/XiBC2aCzGFr8J7nwhazuc3C0A0Ui8JMFeT+ypjTl0tvC
uRSaHikQT30Xa7AQGcENDOxrYSmLTnl9iodARTKH2mqjTfdDqvR94i2wkb2vfVLTtfFDOeUezSPf
b8jLbOyxxc2IfH9dYpf5neNMBb8uJfUGIJ3Ri/4SQpkzoNC3hk+j/CtggZadIiucSYovuztrrhdi
MJGUCwwQBxq1TOx7/j3N9z7WSIcVDOpqtAZFzVPCy9LTQMjs+qgf2gRZcCqb6Lz9ItF5561Zxr/o
bYOjc9mS01G+6UUdBOyQD7dN0q2lkUvOwnDz2kBxHcCiJWSXnO203Pkm0UXQaTVDYKIPFtFF0Qv6
EyErlrAIkUBCxyLdSTm0b6MkN6ISbq/t6jLdEASVMVciGHYZKptwXUqwlSlTnkEvQlSCFGuN/vZC
e7PRQR9fTrRbxvyMPGDSBIC/cKJ7Gy6DQovIvl7VwnJXiIr3EKsaOXDu266cwZumZsaDSFXyXtFh
OXzOdOZp/JHwGcPYs+dE6mg28/H6r0uKta2JxFGlCQq0TGZLCfUTJC54Doa3KPkL/BFeMexZvv3M
HJgTtoXPFvct+LbHPGKoF5erOQ5wsSxBaAYvztVAKdYrFzoI22c//U5PSd+9LqV4RIXW81beErEc
HeDm3iyNuf+UAdQ0ceaqy+1znRK0V+IsBHi0JXwpGmyCmwKDkf+LFiRJBruAkARItpSiNUHJypm/
ZX/MGfKFwhW19uPoys9ez+XpEMWKKVG+E4oWbVRgzBIHmyu3MDvzuHSdOIzXmTb3muzX4fngebFG
k3sD/KGkf1cIYrU3w8WT8Y0iwirLUysvoAPZY0lxgkswepZlkxqmejTd1KXCB2I8oTYpf8Ov8HoX
jMhNKMWVCOmIPPbCs8tv5ijqEhHq12daaEdrJHflMcBTxWSZfSbIWmSn1Q+tB7rWP9sbDzuyaEBE
8EfmS9rfvDT64G7Hbi4EgVVEbIEe8057eSrmYs9wKaahd0qnoer4TkHF4GlIqlittC8obsHxSnA6
I1dGoXLstXlbMUSWKeoq5PxYyvVmvvVYD3vzK9dBXgzjcvF0sXOen5Spd3EjwKLOYs/I22RvK0U0
YcHu7TuVE+QEES1rlcGFcYq35b/+TG4Ix7vQSvKU2Vxcvp5Lse56IKtPkT2KWNNqOo5Jbw5cn+iS
JmaBe4UQlwFcGn+R/uVmxITXzuZEQUpb7TP0T2kLNJpUsqHpWPCvR7805fVMNlCkdHbqZ9GwLqvX
um2NnzzvBkDAOAJGqqCo2j8vW05yHKMdKS28gvDtolkTbJ38EqQDJ6viGEo2EX/QDtyOK3Ctp247
3IodTJi/Ml47U7FC+TeXEA6gdpdn5xn+TE5vqtr8eyeUHUUB0H0kq87uwGeFvH4kZ1OXgfUz4RJR
/pGtMyb/reX6f466LOOUWq8TFLrKd0vMW6V8AikgeQJASB8/++wim01YzxUUj2i62a9lco9RO0lM
50oxt8D7uSVal7YsGXEFBIc9ghz0Vn+Km7spzN3pAyR4u2SnnfEzSaRNgM/vxey/P4lIXtn8kP7P
d0xsPzZ6TrDZXthiAPV+ZBDIl87grU1C8n8URY71lX+Z4SG84NBeOt4vr/hYgkxLLWzrDn/npQwP
uTb+QWzVuc7+9LSomKRE9xEVu4V1Xm+eaqkX8NCNWKAnSCnHyPGNVgeho/FB5ccphkF1ai0+VR/m
mQQubvpMjD7raeyB2sUU/Hcf/OEH4PWPRe7jS9n1mosGN68vGZNr9+r6T/+g1alaDkDfDe3Zt9Zl
AJNtENjcJ5JzFTLmNaGy5UPyWA3ANFpxd7xz0AiAS2mfsbDxqxC7ijvRwzEw2HKYsXeoK9JP9BG2
d/CsNOixK1xV0SS01czIHTH7/cWoTaRh1vTSTcIHx5AelyF5QYW7nA3KRO9bAbiV6ckXnf9IK754
iCGk0Z8aRmxw4XF7GZkX9gkX6iyyf1cyZYJC/lZcnga5vA+nFTbgBYIhr7USXd/6qqA3rEBnh/SZ
nPoieyiyLRbeyN7LklI3w57Q9Y1AbMQNGmDENGy53D6t4xSM54gZeIfbVc5StyzoBSbEI9GGFjMx
Bl2cZN55QAOQlcd2XNH2136wDVAAsl3cdP4wqCFgvSG6O0qqufSq7A31aJqYGXglub9KxiT63Too
6aa0QsmdalWGWWw9UCD1TtgxcVLcAPIA/nfWDm++cchjiMHYtQ8NUPyrXiEAcAenZiQ7K3Ps9iG4
2DZGOWqL8n9fZJFftSfhT6faxgFzNurVVjBYhmr+ap4x7pOcIMUanyM5s9v3eYbIqpXeomT0h1TM
EZqaL3UqUUBl30H3jfq4ZCvZ2yA2BafiaaqVl5Yras4nAHd5apFXFh/g3ZTRRjof0gte6PQSWNbs
8WxwKMAScRa9oRX4wxBGx9U3mri/vmMAgmQfLtKGrmVjDEtRuMo1o067kIqJeHPtHh4EHuW20oT5
+ttGdSeufF7jGNd7/iVQKfNZ7B1vxdK0DlRx14IZWcynxNvrkSMpEF+HZzb3eZZY5B4d2zoIjAL+
dqgXqTght96cngosg8NTwhKLvgQwRRS9WDNuBQNfPq9y23YlsmF3SwtlQ9iLFScT0gFJxN/0JWxT
NJTQRyZWgf0TRYbXb2iTwjbaKDnSUaTEChzV2c4tFapnzzYihWm3i1T5shymqmTLeeWm8qWIWZBq
svd9As3DFc/v4s/2yHXnylyN9MQF8Y5jxrOqCVzSXnUaGnIIROAy4LfgO8gQ8CXrMWtEMuRDcoJa
nY9mNFoTBSCHP75U1w/80odzPUYCOMX4BkfdPGmqvihaXkJmVAsCvXuYjsN4nzi3E3DPbP3u3mNb
T1aEz+3Dwqh7+N2GjuB88hMD+B5SXxvVWhyyIzKG0hUrWECk4uX9YRgtSrpRndQ9c4di3T4VmYYT
SkuYCeM6xoEENJQeqoum0ZoSbLCBaQ3RguuKvzDzsqpcNROrAg81Zh1gxg4PcbABvt9grSApjEPd
4aM7lqWe6WntvayR9GrgVYZaLnFrMdtLhCR2KASgwJy3QTgrPoXu4IpGisW3XDBc/adbZiZJ3vaf
YQyxJMHa80PTM1e/rvCY9oRHj+G0STebTUTw2W2q6XdmWfHBQZ5r5VpGC7FzXTjthU5p5XyVdv+y
n4PX91m4eHRxtOKpedZTPKOKFjvwWCZcf926ASJPaZO0Q3wtTIMij2m3v0JG+XWbojIsWXoOY3Iw
Lne/ca6lH7FU3Y/BAdQWjdnprowiE7+06nwUKfX7evhuJYeh3ynGOAFRCdMhHvSC3A8zfAkRrWvs
EGX0uJ2z+sV8Cdnyb9I3GtsVD68WZZbj/gwlCqMGwde5mDW5ZqJchh7eXNfEX0Mr6sYP3yl5Qnp8
LREe4JUh30uBxG70ulkMCMy+Bb0EzLjNQnOOjHGUjZRiZQwumJqAzJ7Toqg9k8+f0fU7KpF/xL1B
23bVeRz96q8Id8aHJZCwyz0WsRgUwIAUe4r6huvU4BjEwbjKBGz7EWaVIb5oxp/2ilOZo98FM9Uy
CGr3oQ4v8rIFYjoSI1SLWN3lQOhG4aY7zRFC1MZS+ldaOEMxHo0pZ6HI7gvaUgHh5/RrvJfkpuXz
Ta/QV0+282rozDayrcfM75NJtqKzJ8DLt7rgHWrttXOMfERaztrzM1GYwyd6kxEqfcYStIrLYXi+
GD2GQlsamKuvWOcz8SHnjH0TmxOTzvWozzSbGXynsVyQzdylpye+1jV6G6yHppw9m36mxjVwXHr3
RmEqlxFyoSBKq9RTOtTNsHzbIqQE+GObNzkEcjvH0aNS+dFMFJKDguRINKEuz4a8Tt9mjFEHAeTJ
YCB31EcaHurtiQQT79ybrpdfsm4bpnwRrMc1rJIWlSMXOdnb1k8EmBhVBFgJ/1V2LHbM7gnOYiu6
YYpSatY/n6IYEByEJpfMQDliRRPavh+9tawgX3uLG8CaCZyYTUh2WB0vCKIGCPzoN4dxDVaCuj5g
tUE1xEwCyaiksXR8dsnh1WmGGcs2iwbeRw8dodNQ2mOGMNUPmUZXGbmbvJml2HR/KV4sngIn07Y3
x8/Sf0WI5dcAfUzuiVLh10XZPfn9Q06UpFDSFeA1tEPOGYZvoIq4Eqt3Wci7ujUe+ATpoukluwot
C2bZEpXnLMrRM5lBfa5ULtc6VmGJ8yXoLd3ANE3n9XpRFnXWm6cFZyPLBJZIHC3pt21q19JThRnt
nW3oyIbJr7cWfSvAT6qub9pa7pL1Y8J/KJ6sRp6OmnGapFOy1DhJjLYwZJWjDwTXHHnZzDoLKJEM
bebaOhmlTyLihf5aJKssIsFBkm8RbcBKE2NEwlT6e3O7dMPjdTtUlPDKfOB1Nl9dZdzY58Jd1UEa
nu1aN+nKujTyiOQV9w2wyCY1Q8q58/5FEl8rYHD/v/osvAswzSwlzuhLnHhlxW4QmYmbmDCilA8k
UUuXmGhcvNAF/DbfCm5GqSNiF7JntY2XI9ZjSjDGXzptvGba21UufOyft4i/n7g7akCsvtpibrFd
8aIYa7XYEgU2AFn/OWyYjzvlvVQ2tILvZJiYFk2brPMr1Cp1mgpPL5vJfIud7cV9WI4atb/ap/5x
SIIwX7bCF2XrLXzpXrgGVqNI39PPTUGcieUvy5YzrrDFwhZwFtmWHMrBRlOhGc4pgZMGx6CrBRSB
F0/8PrMsy7uHbQNovhFV9ZnKXroFWXz2wxpOx7/oJR2LNwpiStULVXmHy0ImI5xg52aqI4HmVChH
FHxTn32dJrmBZll2BV0xt6wuXt+EiJvvBzY49Q+JvwtGlQLK/tQoT0lFJNioJZVxsHhu4r28oxZy
Wpx7Ngb4hC5lZIoaXIVxNYUxjFVhMDGqT5Z1vRXynP/DRI6M86KxVFz9BLxjqDr2o713Ciz3dXM+
Uk6CBtkZINZ8Sn8XgeWTGNrjJOcS2YAcZh9kyuPiWdfnhpq/A5oismbzjJg6vGgQjN/2p0HfEGqz
F4V5FeZDvd1bIictcnjjiwqobZ2YwaE+XeIAx7TI68YktMvtvtd8G2mBORls62BSzgV5aItplB1T
d0dUNRtragiPK9f8woJ+1eQZVdhVSgVrGhgJYC8XqBWtTcFoGfdGhISS3XR4MtXPq2FH6rxKAjTP
XERgi6HB4j5IothHQx5pEhTefX5+uWfzp6gsS9VyYhI3fj+tX+zib43eALwmT5kZcuU+xP6NEK3k
XLEtf6Ut+VOjHP68rewTnV12vCgVjYJePcuFY0j6KgWPPj/D1GX1zCWJzbKyRUAK
`protect end_protected
